magic
tech sky130A
timestamp 1636366393
<< pwell >>
rect -752 3772 -601 3831
rect -744 3771 -601 3772
rect 308 -775 419 -732
<< nmos >>
rect 56 -298 156 -280
rect 56 -446 156 -428
rect 56 -612 156 -594
rect 54 -765 154 -747
rect 53 -919 153 -901
<< ndiff >>
rect 56 -248 156 -235
rect 56 -266 98 -248
rect 116 -266 156 -248
rect 56 -280 156 -266
rect 56 -312 156 -298
rect 56 -330 98 -312
rect 116 -330 156 -312
rect 56 -343 156 -330
rect 56 -396 156 -383
rect 56 -414 98 -396
rect 116 -414 156 -396
rect 56 -428 156 -414
rect 56 -460 156 -446
rect 56 -478 98 -460
rect 116 -478 156 -460
rect 56 -491 156 -478
rect 56 -562 156 -549
rect 56 -580 98 -562
rect 116 -580 156 -562
rect 56 -594 156 -580
rect 56 -626 156 -612
rect 56 -644 98 -626
rect 116 -644 156 -626
rect 56 -657 156 -644
rect 54 -715 154 -702
rect 54 -733 96 -715
rect 114 -733 154 -715
rect 54 -747 154 -733
rect 54 -779 154 -765
rect 54 -797 96 -779
rect 114 -797 154 -779
rect 54 -810 154 -797
rect 53 -869 153 -856
rect 53 -887 95 -869
rect 113 -887 153 -869
rect 53 -901 153 -887
rect 53 -933 153 -919
rect 53 -951 95 -933
rect 113 -951 153 -933
rect 53 -964 153 -951
<< ndiffc >>
rect 98 -266 116 -248
rect 98 -330 116 -312
rect 98 -414 116 -396
rect 98 -478 116 -460
rect 98 -580 116 -562
rect 98 -644 116 -626
rect 96 -733 114 -715
rect 96 -797 114 -779
rect 95 -887 113 -869
rect 95 -951 113 -933
<< psubdiff >>
rect -752 3810 -601 3831
rect -752 3793 -649 3810
rect -632 3793 -601 3810
rect -752 3772 -601 3793
rect -744 3771 -601 3772
rect 308 -745 419 -732
rect 308 -763 361 -745
rect 379 -763 419 -745
rect 308 -775 419 -763
<< psubdiffcont >>
rect -649 3793 -632 3810
rect 361 -763 379 -745
<< poly >>
rect -3 -280 31 -272
rect -3 -298 5 -280
rect 23 -298 56 -280
rect 156 -298 181 -280
rect -3 -306 31 -298
rect -3 -428 31 -420
rect -3 -446 5 -428
rect 23 -446 56 -428
rect 156 -446 181 -428
rect -3 -454 31 -446
rect -3 -594 31 -586
rect -3 -612 5 -594
rect 23 -612 56 -594
rect 156 -612 181 -594
rect -3 -620 31 -612
rect -5 -747 29 -739
rect -5 -765 3 -747
rect 21 -765 54 -747
rect 154 -765 179 -747
rect -5 -773 29 -765
rect -6 -901 28 -893
rect -6 -919 2 -901
rect 20 -919 53 -901
rect 153 -919 178 -901
rect -6 -927 28 -919
<< polycont >>
rect 5 -298 23 -280
rect 5 -446 23 -428
rect 5 -612 23 -594
rect 3 -765 21 -747
rect 2 -919 20 -901
<< locali >>
rect -4380 4203 -4324 4221
rect -4380 4185 -4362 4203
rect -4344 4185 -4324 4203
rect -4380 4114 -4324 4185
rect -4379 4087 -4324 4114
rect -1824 4188 -1768 4206
rect -1824 4170 -1806 4188
rect -1788 4170 -1768 4188
rect -1824 4099 -1768 4170
rect -4379 4078 -4322 4087
rect -4383 3997 -4322 4078
rect -1823 4072 -1768 4099
rect -1823 4063 -1766 4072
rect -4383 3853 -4320 3997
rect -1827 3982 -1766 4063
rect -4383 3847 -4315 3853
rect -4395 3812 -4312 3847
rect -1827 3812 -1764 3982
rect -4396 3807 -4312 3812
rect -4396 1353 -4309 3807
rect -1807 2650 -1783 3812
rect -766 3811 -599 3842
rect -766 3794 -722 3811
rect -704 3810 -599 3811
rect -704 3794 -649 3810
rect -766 3793 -649 3794
rect -632 3793 -599 3810
rect -766 3766 -599 3793
rect -747 3764 -610 3766
rect 2636 2674 2692 2692
rect 2636 2656 2654 2674
rect 2672 2656 2692 2674
rect -1807 2626 -34 2650
rect -4396 1325 -211 1353
rect -239 -390 -211 1325
rect -58 -180 -34 2626
rect 2636 2585 2692 2656
rect 2637 2558 2692 2585
rect 2637 2549 2694 2558
rect 2633 2380 2694 2549
rect 736 2339 2694 2380
rect -55 -206 -37 -180
rect -153 -231 -37 -206
rect -153 -249 -119 -231
rect -101 -249 -37 -231
rect -153 -281 -37 -249
rect -55 -346 -37 -281
rect -3 -248 300 -240
rect -3 -266 98 -248
rect 116 -266 300 -248
rect -3 -274 300 -266
rect -3 -280 31 -274
rect -3 -298 5 -280
rect 23 -298 31 -280
rect -3 -306 31 -298
rect 90 -312 124 -304
rect 90 -330 98 -312
rect 116 -330 124 -312
rect 90 -346 124 -330
rect -55 -368 124 -346
rect -74 -390 124 -388
rect -239 -396 124 -390
rect -239 -414 98 -396
rect 116 -414 124 -396
rect -239 -418 124 -414
rect -97 -420 124 -418
rect -97 -664 -74 -420
rect -3 -422 124 -420
rect -3 -428 31 -422
rect -3 -446 5 -428
rect 23 -446 31 -428
rect -3 -454 31 -446
rect 90 -460 124 -452
rect 90 -478 98 -460
rect 116 -478 124 -460
rect 90 -495 124 -478
rect 189 -495 209 -274
rect 270 -301 300 -274
rect 270 -346 302 -301
rect 736 -332 777 2339
rect 13729 419 14130 420
rect 13600 414 14130 419
rect 13597 412 14130 414
rect 13529 410 14130 412
rect 13395 390 14130 410
rect 13395 372 13413 390
rect 13431 372 14130 390
rect 13395 355 14130 372
rect 13395 354 13502 355
rect 13538 351 13778 355
rect 90 -527 209 -495
rect 273 -476 302 -346
rect 273 -523 575 -476
rect 544 -525 575 -523
rect 738 -525 777 -332
rect 124 -554 209 -553
rect -3 -560 209 -554
rect -3 -561 291 -560
rect 544 -561 777 -525
rect -3 -562 298 -561
rect -3 -580 98 -562
rect 116 -580 298 -562
rect -3 -588 298 -580
rect -3 -594 31 -588
rect -3 -612 5 -594
rect 23 -612 31 -594
rect -3 -620 31 -612
rect 192 -589 298 -588
rect 90 -626 124 -618
rect 90 -644 98 -626
rect 116 -644 124 -626
rect 90 -664 124 -644
rect -97 -688 124 -664
rect -226 -715 122 -707
rect -226 -733 96 -715
rect 114 -733 122 -715
rect -226 -739 122 -733
rect -226 -981 -194 -739
rect -5 -741 122 -739
rect -5 -747 29 -741
rect -5 -765 3 -747
rect 21 -765 29 -747
rect -5 -773 29 -765
rect 88 -779 122 -771
rect 88 -797 96 -779
rect 114 -797 122 -779
rect 88 -822 122 -797
rect 192 -822 209 -589
rect 248 -636 298 -589
rect 14089 -636 14130 355
rect 248 -677 14130 -636
rect 353 -745 387 -737
rect 353 -763 361 -745
rect 379 -763 387 -745
rect 353 -771 387 -763
rect -134 -861 -46 -838
rect 88 -839 209 -822
rect -134 -863 121 -861
rect -134 -881 -100 -863
rect -82 -869 121 -863
rect -82 -881 95 -869
rect -134 -887 95 -881
rect 113 -887 121 -869
rect -134 -893 121 -887
rect -134 -913 -46 -893
rect -6 -895 121 -893
rect -6 -901 28 -895
rect -6 -919 2 -901
rect 20 -919 28 -901
rect -6 -927 28 -919
rect 87 -933 121 -925
rect 87 -951 95 -933
rect 113 -951 121 -933
rect 87 -977 121 -951
rect -39 -981 420 -977
rect -226 -1013 420 -981
rect -39 -1017 420 -1013
rect -29 -3075 55 -3073
rect -163 -3082 55 -3075
rect 380 -3082 420 -1017
rect -163 -3095 420 -3082
rect -163 -3113 -145 -3095
rect -127 -3113 420 -3095
rect -163 -3122 420 -3113
rect -163 -3130 55 -3122
rect -163 -3131 -56 -3130
rect -20 -3134 55 -3130
<< viali >>
rect -4362 4185 -4344 4203
rect -1806 4170 -1788 4188
rect -722 3794 -704 3811
rect 2654 2656 2672 2674
rect -119 -249 -101 -231
rect 13413 372 13431 390
rect -100 -881 -82 -863
rect -145 -3113 -127 -3095
<< metal1 >>
rect -4380 4207 -4324 4221
rect -4380 4181 -4366 4207
rect -4340 4181 -4324 4207
rect -4380 4143 -4324 4181
rect -1824 4192 -1768 4206
rect -1824 4166 -1810 4192
rect -1784 4166 -1768 4192
rect -1824 4128 -1768 4166
rect -763 3816 -682 3842
rect -763 3789 -726 3816
rect -700 3789 -682 3816
rect -763 3764 -682 3789
rect 2636 2678 2692 2692
rect 2636 2652 2650 2678
rect 2676 2652 2692 2678
rect 2636 2614 2692 2652
rect 13395 394 13473 410
rect 13395 368 13409 394
rect 13435 368 13473 394
rect 13395 354 13473 368
rect -153 -227 -65 -206
rect -153 -253 -123 -227
rect -97 -253 -65 -227
rect -153 -281 -65 -253
rect -134 -859 -46 -838
rect -134 -885 -104 -859
rect -78 -885 -46 -859
rect -134 -913 -46 -885
rect -163 -3091 -85 -3075
rect -163 -3117 -149 -3091
rect -123 -3117 -85 -3091
rect -163 -3131 -85 -3117
<< via1 >>
rect -4366 4203 -4340 4207
rect -4366 4185 -4362 4203
rect -4362 4185 -4344 4203
rect -4344 4185 -4340 4203
rect -4366 4181 -4340 4185
rect -1810 4188 -1784 4192
rect -1810 4170 -1806 4188
rect -1806 4170 -1788 4188
rect -1788 4170 -1784 4188
rect -1810 4166 -1784 4170
rect -726 3811 -700 3816
rect -726 3794 -722 3811
rect -722 3794 -704 3811
rect -704 3794 -700 3811
rect -726 3789 -700 3794
rect 2650 2674 2676 2678
rect 2650 2656 2654 2674
rect 2654 2656 2672 2674
rect 2672 2656 2676 2674
rect 2650 2652 2676 2656
rect 13409 390 13435 394
rect 13409 372 13413 390
rect 13413 372 13431 390
rect 13431 372 13435 390
rect 13409 368 13435 372
rect -123 -231 -97 -227
rect -123 -249 -119 -231
rect -119 -249 -101 -231
rect -101 -249 -97 -231
rect -123 -253 -97 -249
rect -104 -863 -78 -859
rect -104 -881 -100 -863
rect -100 -881 -82 -863
rect -82 -881 -78 -863
rect -104 -885 -78 -881
rect -149 -3095 -123 -3091
rect -149 -3113 -145 -3095
rect -145 -3113 -127 -3095
rect -127 -3113 -123 -3095
rect -149 -3117 -123 -3113
<< metal2 >>
rect -4380 4207 -4324 4221
rect -4380 4181 -4366 4207
rect -4340 4181 -4324 4207
rect -4380 4108 -4324 4181
rect -4380 4079 -4366 4108
rect -4338 4079 -4324 4108
rect -4380 4067 -4324 4079
rect -1824 4192 -1768 4206
rect -1824 4166 -1810 4192
rect -1784 4166 -1768 4192
rect -1824 4093 -1768 4166
rect -1824 4064 -1810 4093
rect -1782 4064 -1768 4093
rect -1824 4052 -1768 4064
rect -763 3816 -682 3842
rect -763 3788 -727 3816
rect -699 3788 -682 3816
rect -763 3764 -682 3788
rect 2636 2678 2692 2692
rect 2636 2652 2650 2678
rect 2676 2652 2692 2678
rect 2636 2579 2692 2652
rect 2636 2550 2650 2579
rect 2678 2550 2692 2579
rect 2636 2538 2692 2550
rect 13395 396 13549 410
rect 13395 394 13508 396
rect 13395 368 13409 394
rect 13435 368 13508 394
rect 13537 368 13549 396
rect 13395 354 13549 368
rect -153 -226 -65 -206
rect -153 -254 -124 -226
rect -96 -254 -65 -226
rect -153 -281 -65 -254
rect -134 -859 -46 -838
rect -134 -885 -104 -859
rect -78 -885 -46 -859
rect -134 -913 -46 -885
rect -110 -1135 -56 -913
rect -110 -1183 1399 -1135
rect -163 -3089 -9 -3075
rect -163 -3091 -50 -3089
rect -163 -3117 -149 -3091
rect -123 -3117 -50 -3091
rect -21 -3117 -9 -3089
rect -163 -3131 -9 -3117
rect 1351 -4539 1399 -1183
rect 1811 -4521 1976 -4472
rect 1811 -4539 1868 -4521
rect 1351 -4587 1868 -4539
rect 1811 -4590 1868 -4587
rect 1936 -4590 1976 -4521
rect 1811 -4649 1976 -4590
<< via2 >>
rect -4366 4079 -4338 4108
rect -1810 4064 -1782 4093
rect -727 3789 -726 3816
rect -726 3789 -700 3816
rect -700 3789 -699 3816
rect -727 3788 -699 3789
rect 2650 2550 2678 2579
rect 13508 368 13537 396
rect -124 -227 -96 -226
rect -124 -253 -123 -227
rect -123 -253 -97 -227
rect -97 -253 -96 -227
rect -124 -254 -96 -253
rect -50 -3117 -21 -3089
rect 1868 -4590 1936 -4521
<< metal3 >>
rect -5523 17055 -4738 17057
rect -5523 17025 -2927 17055
rect -740 17030 -683 17077
rect -5523 17020 -2930 17025
rect -5523 17018 -4738 17020
rect -4804 4110 -3524 14409
rect -4804 4087 -4368 4110
rect -4380 4077 -4368 4087
rect -4336 4087 -3524 4110
rect -4336 4077 -4324 4087
rect -4380 4067 -4324 4077
rect -3944 3827 -3905 4087
rect -3943 -1419 -3905 3827
rect -2969 722 -2930 17020
rect -2186 4095 -906 14399
rect -2186 4077 -1812 4095
rect -1824 4062 -1812 4077
rect -1780 4077 -906 4095
rect -1780 4062 -1768 4077
rect -1824 4052 -1768 4062
rect -1388 3847 -1349 4077
rect -1388 3743 -1347 3847
rect -743 3839 -683 17030
rect -743 3816 -681 3839
rect -743 3788 -727 3816
rect -699 3788 -681 3816
rect -743 3765 -681 3788
rect -744 3743 -681 3765
rect -1388 3736 -681 3743
rect -1388 3686 -685 3736
rect 2304 2605 3584 12927
rect 2424 2604 3436 2605
rect 2578 2581 2763 2604
rect 2578 2556 2648 2581
rect 2636 2548 2648 2556
rect 2680 2556 2763 2581
rect 2680 2548 2692 2556
rect 2636 2538 2692 2548
rect 3071 2307 3106 2604
rect 3070 1277 3106 2307
rect 13808 1277 13844 3144
rect 3070 1241 13844 1277
rect 3010 825 13554 1018
rect 13808 825 13844 1241
rect 3010 789 13844 825
rect -2969 683 -356 722
rect -395 -223 -356 683
rect 3010 398 13554 789
rect 3010 366 13506 398
rect 13539 366 13554 398
rect 3010 184 13554 366
rect -153 -223 -65 -206
rect -395 -226 -65 -223
rect -395 -254 -124 -226
rect -96 -254 -65 -226
rect -395 -262 -65 -254
rect -177 -263 -65 -262
rect -153 -281 -65 -263
rect -133 -282 -92 -281
rect -3943 -1420 760 -1419
rect -3943 -1457 826 -1420
rect 781 -1630 826 -1457
rect 781 -1962 817 -1630
rect 16523 -1962 16559 3105
rect 781 -1998 16559 -1962
rect -10313 -2660 -70 -2466
rect 781 -2660 817 -1998
rect -10313 -2696 817 -2660
rect -10313 -3037 -70 -2696
rect -10313 -3075 -24 -3037
rect -10313 -3087 -9 -3075
rect -10313 -3119 -52 -3087
rect -19 -3119 -9 -3087
rect -10313 -3131 -9 -3119
rect -10313 -3177 -24 -3131
rect -10313 -3290 -70 -3177
rect 1811 -4503 1976 -4472
rect 1811 -4521 2140 -4503
rect 1811 -4590 1868 -4521
rect 1936 -4590 2140 -4521
rect 1811 -4614 2140 -4590
rect 1811 -4649 1976 -4614
<< via3 >>
rect -4368 4108 -4336 4110
rect -4368 4079 -4366 4108
rect -4366 4079 -4338 4108
rect -4338 4079 -4336 4108
rect -4368 4077 -4336 4079
rect -1812 4093 -1780 4095
rect -1812 4064 -1810 4093
rect -1810 4064 -1782 4093
rect -1782 4064 -1780 4093
rect -1812 4062 -1780 4064
rect 2648 2579 2680 2581
rect 2648 2550 2650 2579
rect 2650 2550 2678 2579
rect 2678 2550 2680 2579
rect 2648 2548 2680 2550
rect 13506 396 13539 398
rect 13506 368 13508 396
rect 13508 368 13537 396
rect 13537 368 13539 396
rect 13506 366 13539 368
rect -52 -3089 -19 -3087
rect -52 -3117 -50 -3089
rect -50 -3117 -21 -3089
rect -21 -3117 -19 -3089
rect -52 -3119 -19 -3117
<< mimcap >>
rect -4389 4289 -3889 14244
rect -4389 4256 -4366 4289
rect -4333 4256 -3889 4289
rect -4389 4243 -3889 4256
rect -1833 4274 -1333 14229
rect -1833 4241 -1810 4274
rect -1777 4241 -1333 4274
rect -1833 4228 -1333 4241
rect 2627 2760 3127 12715
rect 2627 2727 2650 2760
rect 2683 2727 3127 2760
rect 2627 2715 3127 2727
rect 3372 401 13372 845
rect 3372 368 13327 401
rect 13360 368 13372 401
rect 3372 345 13372 368
rect -10186 -3084 -186 -2640
rect -10186 -3117 -231 -3084
rect -198 -3117 -186 -3084
rect -10186 -3140 -186 -3117
<< mimcapcontact >>
rect -4366 4256 -4333 4289
rect -1810 4241 -1777 4274
rect 2650 2727 2683 2760
rect 13327 368 13360 401
rect -231 -3117 -198 -3084
<< metal4 >>
rect -4372 4289 -4327 4298
rect -4372 4256 -4366 4289
rect -4333 4256 -4327 4289
rect -4372 4221 -4327 4256
rect -1816 4274 -1771 4283
rect -1816 4241 -1810 4274
rect -1777 4241 -1771 4274
rect -4380 4110 -4324 4221
rect -1816 4206 -1771 4241
rect -4380 4077 -4368 4110
rect -4336 4077 -4324 4110
rect -4380 4068 -4324 4077
rect -1824 4095 -1768 4206
rect -1824 4062 -1812 4095
rect -1780 4062 -1768 4095
rect -1824 4053 -1768 4062
rect 2644 2760 2689 2769
rect 2644 2727 2650 2760
rect 2683 2727 2689 2760
rect 2644 2692 2689 2727
rect 2636 2581 2692 2692
rect 2636 2548 2648 2581
rect 2680 2548 2692 2581
rect 2636 2539 2692 2548
rect 13395 407 13548 410
rect 13318 401 13548 407
rect 13318 368 13327 401
rect 13360 398 13548 401
rect 13360 368 13506 398
rect 13318 366 13506 368
rect 13539 366 13548 398
rect 13318 362 13548 366
rect 13395 354 13548 362
rect -163 -3078 -10 -3075
rect -240 -3084 -10 -3078
rect -240 -3117 -231 -3084
rect -198 -3087 -10 -3084
rect -198 -3117 -52 -3087
rect -240 -3119 -52 -3117
rect -19 -3119 -10 -3087
rect -240 -3123 -10 -3119
rect -163 -3131 -10 -3123
<< labels >>
rlabel metal3 s -139 -241 -139 -241 4 io_analog[2]
rlabel metal3 s -715 3807 -715 3807 4 vssa1
rlabel metal2 s -87 -904 -87 -904 4 vccd1
rlabel metal3 s 800 -1979 800 -1979 4 io_analog[0]
rlabel metal3 s 13823 1255 13823 1255 4 io_analog[1]
<< end >>
