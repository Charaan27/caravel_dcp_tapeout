magic
tech sky130A
timestamp 1636377389
<< metal2 >>
rect 262 -400 318 240
rect 853 -400 909 240
rect 1444 -400 1500 240
rect 2035 -400 2091 240
rect 2626 -400 2682 240
rect 3217 -400 3273 240
rect 3808 -400 3864 240
rect 4399 -400 4455 240
rect 4990 -400 5046 240
rect 5581 -400 5637 240
rect 6172 -400 6228 240
rect 6763 -400 6819 240
rect 7354 -400 7410 240
rect 7945 -400 8001 240
rect 8536 -400 8592 240
rect 9127 -400 9183 240
rect 9718 -400 9774 240
rect 10309 -400 10365 240
rect 10900 -400 10956 240
rect 11491 -400 11547 240
rect 12082 -400 12138 240
rect 12673 -400 12729 240
rect 13264 -400 13320 240
rect 13855 -400 13911 240
rect 14446 -400 14502 240
rect 15037 -400 15093 240
rect 15628 -400 15684 240
rect 16219 -400 16275 240
rect 16810 -400 16866 240
rect 17401 -400 17457 240
rect 17992 -400 18048 240
rect 18583 -400 18639 240
rect 19174 -400 19230 240
rect 19765 -400 19821 240
rect 20356 -400 20412 240
rect 20947 -400 21003 240
rect 21538 -400 21594 240
rect 22129 -400 22185 240
rect 22720 -400 22776 240
rect 23311 -400 23367 240
rect 23902 -400 23958 240
rect 24493 -400 24549 240
rect 25084 -400 25140 240
rect 25675 -400 25731 240
rect 26266 -400 26322 240
rect 26857 -400 26913 240
rect 27448 -400 27504 240
rect 28039 -400 28095 240
rect 28630 -400 28686 240
rect 29221 -400 29277 240
rect 29812 -400 29868 240
rect 30403 -400 30459 240
rect 30994 -400 31050 240
rect 31585 -400 31641 240
rect 32176 -400 32232 240
rect 32767 -400 32823 240
rect 33358 -400 33414 240
rect 33949 -400 34005 240
rect 34540 -400 34596 240
rect 35131 -400 35187 240
rect 35722 -400 35778 240
rect 36313 -400 36369 240
rect 36904 -400 36960 240
rect 37495 -400 37551 240
rect 38086 -400 38142 240
rect 38677 -400 38733 240
rect 39268 -400 39324 240
rect 39859 -400 39915 240
rect 40450 -400 40506 240
rect 41041 -400 41097 240
rect 41632 -400 41688 240
rect 42223 -400 42279 240
rect 42814 -400 42870 240
rect 43405 -400 43461 240
rect 43996 -400 44052 240
rect 44587 -400 44643 240
rect 45178 -400 45234 240
rect 45769 -400 45825 240
rect 46360 -400 46416 240
rect 46951 -400 47007 240
rect 47542 -400 47598 240
rect 48133 -400 48189 240
rect 48724 -400 48780 240
rect 49315 -400 49371 240
rect 49906 -400 49962 240
rect 50497 -400 50553 240
rect 51088 -400 51144 240
rect 51679 -400 51735 240
rect 52270 -400 52326 240
rect 52861 -400 52917 240
rect 53452 -400 53508 240
rect 54043 -400 54099 240
rect 54634 -400 54690 240
rect 55225 -400 55281 240
rect 55816 -400 55872 240
rect 56407 -400 56463 240
rect 56998 -400 57054 240
rect 57589 -400 57645 240
rect 58180 -400 58236 240
rect 58771 -400 58827 240
rect 59362 -400 59418 240
rect 59953 -400 60009 240
rect 60544 -400 60600 240
rect 61135 -400 61191 240
rect 61726 -400 61782 240
rect 62317 -400 62373 240
rect 62908 -400 62964 240
rect 63499 -400 63555 240
rect 64090 -400 64146 240
rect 64681 -400 64737 240
rect 65272 -400 65328 240
rect 65863 -400 65919 240
rect 66454 -400 66510 240
rect 67045 -400 67101 240
rect 67636 -400 67692 240
rect 68227 -400 68283 240
rect 68818 -400 68874 240
rect 69409 -400 69465 240
rect 70000 -400 70056 240
rect 70591 -400 70647 240
rect 71182 -400 71238 240
rect 71773 -400 71829 240
rect 72364 -400 72420 240
rect 72955 -400 73011 240
rect 73546 -400 73602 240
rect 74137 -400 74193 240
rect 74728 -400 74784 240
rect 75319 -400 75375 240
rect 75910 -400 75966 240
rect 76501 -400 76557 240
rect 77092 -400 77148 240
rect 77683 -400 77739 240
rect 78274 -400 78330 240
rect 78865 -400 78921 240
rect 79456 -400 79512 240
rect 80047 -400 80103 240
rect 80638 -400 80694 240
rect 81229 -400 81285 240
rect 81820 -400 81876 240
rect 82411 -400 82467 240
rect 83002 -400 83058 240
rect 83593 -400 83649 240
rect 84184 -400 84240 240
rect 84775 -400 84831 240
rect 85366 -400 85422 240
rect 85957 -400 86013 240
rect 86548 -400 86604 240
rect 87139 -400 87195 240
rect 87730 -400 87786 240
rect 88321 -400 88377 240
rect 88912 -400 88968 240
rect 89503 -400 89559 240
rect 90094 -400 90150 240
rect 90685 -400 90741 240
rect 91276 -400 91332 240
rect 91867 -400 91923 240
rect 92458 -400 92514 240
rect 93049 -400 93105 240
rect 93640 -400 93696 240
rect 94231 -400 94287 240
rect 94822 -400 94878 240
rect 95413 -400 95469 240
rect 96004 -400 96060 240
rect 96595 -400 96651 240
rect 97186 -400 97242 240
rect 97777 -400 97833 240
rect 98368 -400 98424 240
rect 98959 -400 99015 240
rect 99550 -400 99606 240
rect 100141 -400 100197 240
rect 100732 -400 100788 240
rect 101323 -400 101379 240
rect 101914 -400 101970 240
rect 102505 -400 102561 240
rect 103096 -400 103152 240
rect 103687 -400 103743 240
rect 104278 -400 104334 240
rect 104869 -400 104925 240
rect 105460 -400 105516 240
rect 106051 -400 106107 240
rect 106642 -400 106698 240
rect 107233 -400 107289 240
rect 107824 -400 107880 240
rect 108415 -400 108471 240
rect 109006 -400 109062 240
rect 109597 -400 109653 240
rect 110188 -400 110244 240
rect 110779 -400 110835 240
rect 111370 -400 111426 240
rect 111961 -400 112017 240
rect 112552 -400 112608 240
rect 113143 -400 113199 240
rect 113734 -400 113790 240
rect 114325 -400 114381 240
rect 114916 -400 114972 240
rect 115507 -400 115563 240
rect 116098 -400 116154 240
rect 116689 -400 116745 240
rect 117280 -400 117336 240
rect 117871 -400 117927 240
rect 118462 -400 118518 240
rect 119053 -400 119109 240
rect 119644 -400 119700 240
rect 120235 -400 120291 240
rect 120826 -400 120882 240
rect 121417 -400 121473 240
rect 122008 -400 122064 240
rect 122599 -400 122655 240
rect 123190 -400 123246 240
rect 123781 -400 123837 240
rect 124372 -400 124428 240
rect 124963 -400 125019 240
rect 125554 -400 125610 240
rect 126145 -400 126201 240
rect 126736 -400 126792 240
rect 127327 -400 127383 240
rect 127918 -400 127974 240
rect 128509 -400 128565 240
rect 129100 -400 129156 240
rect 129691 -400 129747 240
rect 130282 -400 130338 240
rect 130873 -400 130929 240
rect 131464 -400 131520 240
rect 132055 -400 132111 240
rect 132646 -400 132702 240
rect 133237 -400 133293 240
rect 133828 -400 133884 240
rect 134419 -400 134475 240
rect 135010 -400 135066 240
rect 135601 -400 135657 240
rect 136192 -400 136248 240
rect 136783 -400 136839 240
rect 137374 -400 137430 240
rect 137965 -400 138021 240
rect 138556 -400 138612 240
rect 139147 -400 139203 240
rect 139738 -400 139794 240
rect 140329 -400 140385 240
rect 140920 -400 140976 240
rect 141511 -400 141567 240
rect 142102 -400 142158 240
rect 142693 -400 142749 240
rect 143284 -400 143340 240
rect 143875 -400 143931 240
rect 144466 -400 144522 240
rect 145057 -400 145113 240
rect 145648 -400 145704 240
rect 146239 -400 146295 240
rect 146830 -400 146886 240
rect 147421 -400 147477 240
rect 148012 -400 148068 240
rect 148603 -400 148659 240
rect 149194 -400 149250 240
rect 149785 -400 149841 240
rect 150376 -400 150432 240
rect 150967 -400 151023 240
rect 151558 -400 151614 240
rect 152149 -400 152205 240
rect 152740 -400 152796 240
rect 153331 -400 153387 240
rect 153922 -400 153978 240
rect 154513 -400 154569 240
rect 155104 -400 155160 240
rect 155695 -400 155751 240
rect 156286 -400 156342 240
rect 156877 -400 156933 240
rect 157468 -400 157524 240
rect 158059 -400 158115 240
rect 158650 -400 158706 240
rect 159241 -400 159297 240
rect 159832 -400 159888 240
rect 160423 -400 160479 240
rect 161014 -400 161070 240
rect 161605 -400 161661 240
rect 162196 -400 162252 240
rect 162787 -400 162843 240
rect 163378 -400 163434 240
rect 163969 -400 164025 240
rect 164560 -400 164616 240
rect 165151 -400 165207 240
rect 165742 -400 165798 240
rect 166333 -400 166389 240
rect 166924 -400 166980 240
rect 167515 -400 167571 240
rect 168106 -400 168162 240
rect 168697 -400 168753 240
rect 169288 -400 169344 240
rect 169879 -400 169935 240
rect 170470 -400 170526 240
rect 171061 -400 171117 240
rect 171652 -400 171708 240
rect 172243 -400 172299 240
rect 172834 -400 172890 240
rect 173425 -400 173481 240
rect 174016 -400 174072 240
rect 174607 -400 174663 240
rect 175198 -400 175254 240
rect 175789 -400 175845 240
rect 176380 -400 176436 240
rect 176971 -400 177027 240
rect 177562 -400 177618 240
rect 178153 -400 178209 240
rect 178744 -400 178800 240
rect 179335 -400 179391 240
rect 179926 -400 179982 240
rect 180517 -400 180573 240
rect 181108 -400 181164 240
rect 181699 -400 181755 240
rect 182290 -400 182346 240
rect 182881 -400 182937 240
rect 183472 -400 183528 240
rect 184063 -400 184119 240
rect 184654 -400 184710 240
rect 185245 -400 185301 240
rect 185836 -400 185892 240
rect 186427 -400 186483 240
rect 187018 -400 187074 240
rect 187609 -400 187665 240
rect 188200 -400 188256 240
rect 188791 -400 188847 240
rect 189382 -400 189438 240
rect 189973 -400 190029 240
rect 190564 -400 190620 240
rect 191155 -400 191211 240
rect 191746 -400 191802 240
rect 192337 -400 192393 240
rect 192928 -400 192984 240
rect 193519 -400 193575 240
rect 194110 -400 194166 240
rect 194701 -400 194757 240
rect 195292 -400 195348 240
rect 195883 -400 195939 240
rect 196474 -400 196530 240
rect 197065 -400 197121 240
rect 197656 -400 197712 240
rect 198247 -400 198303 240
rect 198838 -400 198894 240
rect 199429 -400 199485 240
rect 200020 -400 200076 240
rect 200611 -400 200667 240
rect 201202 -400 201258 240
rect 201793 -400 201849 240
rect 202384 -400 202440 240
rect 202975 -400 203031 240
rect 203566 -400 203622 240
rect 204157 -400 204213 240
rect 204748 -400 204804 240
rect 205339 -400 205395 240
rect 205930 -400 205986 240
rect 206521 -400 206577 240
rect 207112 -400 207168 240
rect 207703 -400 207759 240
rect 208294 -400 208350 240
rect 208885 -400 208941 240
rect 209476 -400 209532 240
rect 210067 -400 210123 240
rect 210658 -400 210714 240
rect 211249 -400 211305 240
rect 211840 -400 211896 240
rect 212431 -400 212487 240
rect 213022 -400 213078 240
rect 213613 -400 213669 240
rect 214204 -400 214260 240
rect 214795 -400 214851 240
rect 215386 -400 215442 240
rect 215977 -400 216033 240
rect 216568 -400 216624 240
rect 217159 -400 217215 240
rect 217750 -400 217806 240
rect 218341 -400 218397 240
rect 218932 -400 218988 240
rect 219523 -400 219579 240
rect 220114 -400 220170 240
rect 220705 -400 220761 240
rect 221296 -400 221352 240
rect 221887 -400 221943 240
rect 222478 -400 222534 240
rect 223069 -400 223125 240
rect 223660 -400 223716 240
rect 224251 -400 224307 240
rect 224842 -400 224898 240
rect 225433 -400 225489 240
rect 226024 -400 226080 240
rect 226615 -400 226671 240
rect 227206 -400 227262 240
rect 227797 -400 227853 240
rect 228388 -400 228444 240
rect 228979 -400 229035 240
rect 229570 -400 229626 240
rect 230161 -400 230217 240
rect 230752 -400 230808 240
rect 231343 -400 231399 240
rect 231934 -400 231990 240
rect 232525 -400 232581 240
rect 233116 -400 233172 240
rect 233707 -400 233763 240
rect 234298 -400 234354 240
rect 234889 -400 234945 240
rect 235480 -400 235536 240
rect 236071 -400 236127 240
rect 236662 -400 236718 240
rect 237253 -400 237309 240
rect 237844 -400 237900 240
rect 238435 -400 238491 240
rect 239026 -400 239082 240
rect 239617 -400 239673 240
rect 240208 -400 240264 240
rect 240799 -400 240855 240
rect 241390 -400 241446 240
rect 241981 -400 242037 240
rect 242572 -400 242628 240
rect 243163 -400 243219 240
rect 243754 -400 243810 240
rect 244345 -400 244401 240
rect 244936 -400 244992 240
rect 245527 -400 245583 240
rect 246118 -400 246174 240
rect 246709 -400 246765 240
rect 247300 -400 247356 240
rect 247891 -400 247947 240
rect 248482 -400 248538 240
rect 249073 -400 249129 240
rect 249664 -400 249720 240
rect 250255 -400 250311 240
rect 250846 -400 250902 240
rect 251437 -400 251493 240
rect 252028 -400 252084 240
rect 252619 -400 252675 240
rect 253210 -400 253266 240
rect 253801 -400 253857 240
rect 254392 -400 254448 240
rect 254983 -400 255039 240
rect 255574 -400 255630 240
rect 256165 -400 256221 240
rect 256756 -400 256812 240
rect 257347 -400 257403 240
rect 257938 -400 257994 240
rect 258529 -400 258585 240
rect 259120 -400 259176 240
rect 259711 -400 259767 240
rect 260302 -400 260358 240
rect 260893 -400 260949 240
rect 261484 -400 261540 240
rect 262075 -400 262131 240
rect 262666 -400 262722 240
rect 263257 -400 263313 240
rect 263848 -400 263904 240
rect 264439 -400 264495 240
rect 265030 -400 265086 240
rect 265621 -400 265677 240
rect 266212 -400 266268 240
rect 266803 -400 266859 240
rect 267394 -400 267450 240
rect 267985 -400 268041 240
rect 268576 -400 268632 240
rect 269167 -400 269223 240
rect 269758 -400 269814 240
rect 270349 -400 270405 240
rect 270940 -400 270996 240
rect 271531 -400 271587 240
rect 272122 -400 272178 240
rect 272713 -400 272769 240
rect 273304 -400 273360 240
rect 273895 -400 273951 240
rect 274486 -400 274542 240
rect 275077 -400 275133 240
rect 275668 -400 275724 240
rect 276259 -400 276315 240
rect 276850 -400 276906 240
rect 277441 -400 277497 240
rect 278032 -400 278088 240
rect 278623 -400 278679 240
rect 279214 -400 279270 240
rect 279805 -400 279861 240
rect 280396 -400 280452 240
rect 280987 -400 281043 240
rect 281578 -400 281634 240
rect 282169 -400 282225 240
rect 282760 -400 282816 240
rect 283351 -400 283407 240
rect 283942 -400 283998 240
rect 284533 -400 284589 240
rect 285124 -400 285180 240
rect 285715 -400 285771 240
rect 286306 -400 286362 240
rect 286897 -400 286953 240
rect 287488 -400 287544 240
rect 288079 -400 288135 240
rect 288670 -400 288726 240
rect 289261 -400 289317 240
rect 289852 -400 289908 240
rect 290443 -400 290499 240
rect 291034 -400 291090 240
rect 291625 -400 291681 240
<< metal3 >>
rect 8097 351150 10597 352400
rect 34097 351150 36597 352400
rect 60097 351150 62597 352400
rect 82797 351150 85297 352400
rect 85447 351150 86547 352400
rect 86697 351150 87797 352400
rect 87947 351150 90447 352400
rect 108647 351150 111147 352400
rect 111297 351150 112397 352400
rect 112547 351150 113647 352400
rect 113797 351150 116297 352400
rect 159497 351150 161997 352400
rect 162147 351150 163247 352400
rect 163397 351150 164497 352400
rect 164647 351150 167147 352400
rect 206697 351150 209197 352400
rect 232697 351150 235197 352400
rect 255297 351170 257697 352400
rect 260297 351170 262697 352400
rect -400 340121 850 342621
rect 234284 335214 234334 351150
rect 261819 350235 261954 351170
rect 283297 351150 285797 352400
rect 261819 350226 266247 350235
rect 268223 350226 268290 350227
rect 261819 350103 268290 350226
rect 283968 350182 284029 351150
rect 283393 350178 284029 350182
rect 261819 350101 266247 350103
rect 261819 350097 261954 350101
rect 268223 336613 268290 350103
rect 282760 350139 284029 350178
rect 282760 350135 283394 350139
rect 282760 348111 282806 350135
rect 283968 350134 284029 350139
rect 282758 344698 282807 348111
rect 268220 336612 268290 336613
rect 268220 335223 268274 336612
rect 282763 335229 282800 344698
rect 285483 339566 285527 339567
rect 291150 339566 292400 341492
rect 285474 339467 292400 339566
rect 285483 335246 285527 339467
rect 291150 338992 292400 339467
rect 234284 335209 256861 335214
rect 234284 335203 258744 335209
rect 268220 335206 268269 335223
rect 234284 335167 263435 335203
rect -400 321921 830 324321
rect 282760 321277 282800 335229
rect 285481 335223 285530 335246
rect 285481 321251 285532 335223
rect 285483 321228 285532 321251
rect 291170 319892 292400 322292
rect -400 316921 830 319321
rect 291170 314892 292400 317292
rect 291872 313645 292018 314892
rect 290627 313641 292018 313645
rect 271062 313638 285603 313641
rect 290627 313638 292022 313641
rect 271062 313532 292022 313638
rect 271062 313531 285603 313532
rect 290627 313519 292022 313532
rect 291789 313513 292022 313519
rect 291872 313509 292018 313513
rect 291760 294736 292400 294792
rect 291760 294145 292400 294201
rect 291760 293554 292400 293610
rect 291760 292963 292400 293019
rect 291760 292372 292400 292428
rect 291760 291781 292400 291837
rect -400 279721 830 282121
rect -400 274721 830 277121
rect 291170 275281 292400 277681
rect 291170 270281 292400 272681
rect -400 255765 240 255821
rect -400 255174 240 255230
rect -400 254583 240 254639
rect -400 253992 240 254048
rect -400 253401 240 253457
rect -400 252810 240 252866
rect 291760 250025 292400 250081
rect 291760 249434 292400 249490
rect 291760 248843 292400 248899
rect 291760 248252 292400 248308
rect 291760 247661 292400 247717
rect 291760 247070 292400 247126
rect -400 234154 240 234210
rect -400 233563 240 233619
rect -400 232972 240 233028
rect -400 232381 240 232437
rect -400 231790 240 231846
rect -400 231199 240 231255
rect 291760 227814 292400 227870
rect 291760 227223 292400 227279
rect 291760 226632 292400 226688
rect 291760 226041 292400 226097
rect 291760 225450 292400 225506
rect 291760 224859 292400 224915
rect -400 212543 240 212599
rect -400 211952 240 212008
rect -400 211361 240 211417
rect -400 210770 240 210826
rect -400 210179 240 210235
rect -400 209588 240 209644
rect 291760 205603 292400 205659
rect 291760 205012 292400 205068
rect 291760 204421 292400 204477
rect 291760 203830 292400 203886
rect 291760 203239 292400 203295
rect 291760 202648 292400 202704
rect -400 190932 240 190988
rect -400 190341 240 190397
rect -400 189750 240 189806
rect -400 189159 240 189215
rect -400 188568 240 188624
rect -400 187977 240 188033
rect 291760 182392 292400 182448
rect 291760 181801 292400 181857
rect 291760 181210 292400 181266
rect 291760 180619 292400 180675
rect 291760 180028 292400 180084
rect 291760 179437 292400 179493
rect -400 169321 240 169377
rect -400 168730 240 168786
rect -400 168139 240 168195
rect -400 167548 240 167604
rect -400 166957 240 167013
rect -400 166366 240 166422
rect 291760 159781 292400 159837
rect 291760 159190 292400 159246
rect 291760 158599 292400 158655
rect 291760 158008 292400 158064
rect 291760 157417 292400 157473
rect 291760 156826 292400 156882
rect -400 147710 240 147766
rect -400 147119 240 147175
rect -400 146528 240 146584
rect -400 145937 240 145993
rect -400 145346 240 145402
rect -400 144755 240 144811
rect 291760 137570 292400 137626
rect 291760 136979 292400 137035
rect 291760 136388 292400 136444
rect 291760 135797 292400 135853
rect 291760 135206 292400 135262
rect 291760 134615 292400 134671
rect -400 126199 240 126255
rect -400 125608 240 125664
rect -400 125017 240 125073
rect -400 124426 240 124482
rect -400 123835 240 123891
rect -400 123244 240 123300
rect 291170 117615 292400 120015
rect 291170 112615 292400 115015
rect -400 107444 830 109844
rect -400 102444 830 104844
rect 291170 95715 292400 98115
rect 291170 90715 292400 93115
rect -400 86444 830 88844
rect -400 81444 830 83844
rect 291170 73415 292400 75815
rect 291170 68415 292400 70815
rect -400 62388 240 62444
rect -400 61797 240 61853
rect -400 61206 240 61262
rect -400 60615 240 60671
rect -400 60024 240 60080
rect -400 59433 240 59489
rect 291760 47559 292400 47615
rect 291760 46968 292400 47024
rect 291760 46377 292400 46433
rect 291760 45786 292400 45842
rect -400 40777 240 40833
rect -400 40186 240 40242
rect -400 39595 240 39651
rect -400 39004 240 39060
rect -400 38413 240 38469
rect -400 37822 240 37878
rect 291760 25230 292400 25286
rect 291760 24639 292400 24695
rect 291760 24048 292400 24104
rect 291760 23457 292400 23513
rect -400 19166 240 19222
rect -400 18575 240 18631
rect -400 17984 240 18040
rect -400 17393 240 17449
rect -400 16802 240 16858
rect -400 16211 240 16267
rect 291760 12001 292400 12057
rect 291760 11410 292400 11466
rect 291760 10819 292400 10875
rect 291760 10228 292400 10284
rect 291760 9637 292400 9693
rect 291760 9046 292400 9102
rect -400 8455 240 8511
rect 291760 8455 292400 8511
rect -400 7864 240 7920
rect 291760 7864 292400 7920
rect -400 7273 240 7329
rect 291760 7273 292400 7329
rect -400 6682 240 6738
rect 291760 6682 292400 6738
rect -400 6091 240 6147
rect 291760 6091 292400 6147
rect -400 5500 240 5556
rect 291760 5500 292400 5556
rect -400 4909 240 4965
rect 291760 4909 292400 4965
rect -400 4318 240 4374
rect 291760 4318 292400 4374
rect -400 3727 240 3783
rect 291760 3727 292400 3783
rect -400 3136 240 3192
rect 291760 3136 292400 3192
rect -400 2545 240 2601
rect 291760 2545 292400 2601
rect -400 1954 240 2010
rect 291760 1954 292400 2010
rect -400 1363 240 1419
rect 291760 1363 292400 1419
rect -400 772 240 828
rect 291760 772 292400 828
use dcp_tapeout  dcp_tapeout_0
timestamp 1636377260
transform 1 0 268958 0 1 318146
box -10313 -4649 16559 17077
<< labels >>
flabel metal3 s 291760 134615 292400 134671 0 FreeSans 6507 0 0 0 gpio_analog[0]
flabel metal3 s -400 190932 240 190988 0 FreeSans 6507 0 0 0 gpio_analog[10]
flabel metal3 s -400 169321 240 169377 0 FreeSans 6507 0 0 0 gpio_analog[11]
flabel metal3 s -400 147710 240 147766 0 FreeSans 6507 0 0 0 gpio_analog[12]
flabel metal3 s -400 126199 240 126255 0 FreeSans 6507 0 0 0 gpio_analog[13]
flabel metal3 s -400 62388 240 62444 0 FreeSans 6507 0 0 0 gpio_analog[14]
flabel metal3 s -400 40777 240 40833 0 FreeSans 6507 0 0 0 gpio_analog[15]
flabel metal3 s -400 19166 240 19222 0 FreeSans 6507 0 0 0 gpio_analog[16]
flabel metal3 s -400 8455 240 8511 0 FreeSans 6507 0 0 0 gpio_analog[17]
flabel metal3 s 291760 156826 292400 156882 0 FreeSans 6507 0 0 0 gpio_analog[1]
flabel metal3 s 291760 179437 292400 179493 0 FreeSans 6507 0 0 0 gpio_analog[2]
flabel metal3 s 291760 202648 292400 202704 0 FreeSans 6507 0 0 0 gpio_analog[3]
flabel metal3 s 291760 224859 292400 224915 0 FreeSans 6507 0 0 0 gpio_analog[4]
flabel metal3 s 291760 247070 292400 247126 0 FreeSans 6507 0 0 0 gpio_analog[5]
flabel metal3 s 291760 291781 292400 291837 0 FreeSans 6507 0 0 0 gpio_analog[6]
flabel metal3 s -400 255765 240 255821 0 FreeSans 6507 0 0 0 gpio_analog[7]
flabel metal3 s -400 234154 240 234210 0 FreeSans 6507 0 0 0 gpio_analog[8]
flabel metal3 s -400 212543 240 212599 0 FreeSans 6507 0 0 0 gpio_analog[9]
flabel metal3 s 291760 135206 292400 135262 0 FreeSans 6507 0 0 0 gpio_noesd[0]
flabel metal3 s -400 190341 240 190397 0 FreeSans 6507 0 0 0 gpio_noesd[10]
flabel metal3 s -400 168730 240 168786 0 FreeSans 6507 0 0 0 gpio_noesd[11]
flabel metal3 s -400 147119 240 147175 0 FreeSans 6507 0 0 0 gpio_noesd[12]
flabel metal3 s -400 125608 240 125664 0 FreeSans 6507 0 0 0 gpio_noesd[13]
flabel metal3 s -400 61797 240 61853 0 FreeSans 6507 0 0 0 gpio_noesd[14]
flabel metal3 s -400 40186 240 40242 0 FreeSans 6507 0 0 0 gpio_noesd[15]
flabel metal3 s -400 18575 240 18631 0 FreeSans 6507 0 0 0 gpio_noesd[16]
flabel metal3 s -400 7864 240 7920 0 FreeSans 6507 0 0 0 gpio_noesd[17]
flabel metal3 s 291760 157417 292400 157473 0 FreeSans 6507 0 0 0 gpio_noesd[1]
flabel metal3 s 291760 180028 292400 180084 0 FreeSans 6507 0 0 0 gpio_noesd[2]
flabel metal3 s 291760 203239 292400 203295 0 FreeSans 6507 0 0 0 gpio_noesd[3]
flabel metal3 s 291760 225450 292400 225506 0 FreeSans 6507 0 0 0 gpio_noesd[4]
flabel metal3 s 291760 247661 292400 247717 0 FreeSans 6507 0 0 0 gpio_noesd[5]
flabel metal3 s 291760 292372 292400 292428 0 FreeSans 6507 0 0 0 gpio_noesd[6]
flabel metal3 s -400 255174 240 255230 0 FreeSans 6507 0 0 0 gpio_noesd[7]
flabel metal3 s -400 233563 240 233619 0 FreeSans 6507 0 0 0 gpio_noesd[8]
flabel metal3 s -400 211952 240 212008 0 FreeSans 6507 0 0 0 gpio_noesd[9]
flabel metal3 s 291150 338992 292400 341492 0 FreeSans 6507 0 0 0 io_analog[0]
flabel metal3 s 0 340121 850 342621 0 FreeSans 6507 0 0 0 io_analog[10]
flabel metal3 s 283297 351150 285797 352400 0 FreeSans 11166 180 0 0 io_analog[1]
flabel metal3 s 232697 351150 235197 352400 0 FreeSans 11166 180 0 0 io_analog[2]
flabel metal3 s 206697 351150 209197 352400 0 FreeSans 11166 180 0 0 io_analog[3]
flabel metal3 s 164647 351150 167147 352400 0 FreeSans 11166 180 0 0 io_analog[4]
flabel metal3 s 113797 351150 116297 352400 0 FreeSans 11166 180 0 0 io_analog[5]
flabel metal3 s 87947 351150 90447 352400 0 FreeSans 11166 180 0 0 io_analog[6]
flabel metal3 s 60097 351150 62597 352400 0 FreeSans 11166 180 0 0 io_analog[7]
flabel metal3 s 34097 351150 36597 352400 0 FreeSans 11166 180 0 0 io_analog[8]
flabel metal3 s 8097 351150 10597 352400 0 FreeSans 11166 180 0 0 io_analog[9]
flabel metal3 s 159497 351150 161997 352400 0 FreeSans 11166 180 0 0 io_analog[4]
flabel metal3 s 108647 351150 111147 352400 0 FreeSans 11166 180 0 0 io_analog[5]
flabel metal3 s 82797 351150 85297 352400 0 FreeSans 11166 180 0 0 io_analog[6]
flabel metal3 s 163397 351150 164497 352400 0 FreeSans 11166 180 0 0 io_clamp_high[0]
flabel metal3 s 112547 351150 113647 352400 0 FreeSans 11166 180 0 0 io_clamp_high[1]
flabel metal3 s 86697 351150 87797 352400 0 FreeSans 11166 180 0 0 io_clamp_high[2]
flabel metal3 s 162147 351150 163247 352400 0 FreeSans 11166 180 0 0 io_clamp_low[0]
flabel metal3 s 111297 351150 112397 352400 0 FreeSans 11166 180 0 0 io_clamp_low[1]
flabel metal3 s 85447 351150 86547 352400 0 FreeSans 11166 180 0 0 io_clamp_low[2]
flabel metal3 s 291760 1363 292400 1419 0 FreeSans 6507 0 0 0 io_in[0]
flabel metal3 s 291760 204421 292400 204477 0 FreeSans 6507 0 0 0 io_in[10]
flabel metal3 s 291760 226632 292400 226688 0 FreeSans 6507 0 0 0 io_in[11]
flabel metal3 s 291760 248843 292400 248899 0 FreeSans 6507 0 0 0 io_in[12]
flabel metal3 s 291760 293554 292400 293610 0 FreeSans 6507 0 0 0 io_in[13]
flabel metal3 s -400 253992 240 254048 0 FreeSans 6507 0 0 0 io_in[14]
flabel metal3 s -400 232381 240 232437 0 FreeSans 6507 0 0 0 io_in[15]
flabel metal3 s -400 210770 240 210826 0 FreeSans 6507 0 0 0 io_in[16]
flabel metal3 s -400 189159 240 189215 0 FreeSans 6507 0 0 0 io_in[17]
flabel metal3 s -400 167548 240 167604 0 FreeSans 6507 0 0 0 io_in[18]
flabel metal3 s -400 145937 240 145993 0 FreeSans 6507 0 0 0 io_in[19]
flabel metal3 s 291760 3727 292400 3783 0 FreeSans 6507 0 0 0 io_in[1]
flabel metal3 s -400 124426 240 124482 0 FreeSans 6507 0 0 0 io_in[20]
flabel metal3 s -400 60615 240 60671 0 FreeSans 6507 0 0 0 io_in[21]
flabel metal3 s -400 39004 240 39060 0 FreeSans 6507 0 0 0 io_in[22]
flabel metal3 s -400 17393 240 17449 0 FreeSans 6507 0 0 0 io_in[23]
flabel metal3 s -400 6682 240 6738 0 FreeSans 6507 0 0 0 io_in[24]
flabel metal3 s -400 4318 240 4374 0 FreeSans 6507 0 0 0 io_in[25]
flabel metal3 s -400 1954 240 2010 0 FreeSans 6507 0 0 0 io_in[26]
flabel metal3 s 291760 6091 292400 6147 0 FreeSans 6507 0 0 0 io_in[2]
flabel metal3 s 291760 8455 292400 8511 0 FreeSans 6507 0 0 0 io_in[3]
flabel metal3 s 291760 10819 292400 10875 0 FreeSans 6507 0 0 0 io_in[4]
flabel metal3 s 291760 24048 292400 24104 0 FreeSans 6507 0 0 0 io_in[5]
flabel metal3 s 291760 46377 292400 46433 0 FreeSans 6507 0 0 0 io_in[6]
flabel metal3 s 291760 136388 292400 136444 0 FreeSans 6507 0 0 0 io_in[7]
flabel metal3 s 291760 158599 292400 158655 0 FreeSans 6507 0 0 0 io_in[8]
flabel metal3 s 291760 181210 292400 181266 0 FreeSans 6507 0 0 0 io_in[9]
flabel metal3 s 291760 772 292400 828 0 FreeSans 6507 0 0 0 io_in_3v3[0]
flabel metal3 s 291760 203830 292400 203886 0 FreeSans 6507 0 0 0 io_in_3v3[10]
flabel metal3 s 291760 226041 292400 226097 0 FreeSans 6507 0 0 0 io_in_3v3[11]
flabel metal3 s 291760 248252 292400 248308 0 FreeSans 6507 0 0 0 io_in_3v3[12]
flabel metal3 s 291760 292963 292400 293019 0 FreeSans 6507 0 0 0 io_in_3v3[13]
flabel metal3 s -400 254583 240 254639 0 FreeSans 6507 0 0 0 io_in_3v3[14]
flabel metal3 s -400 232972 240 233028 0 FreeSans 6507 0 0 0 io_in_3v3[15]
flabel metal3 s -400 211361 240 211417 0 FreeSans 6507 0 0 0 io_in_3v3[16]
flabel metal3 s -400 189750 240 189806 0 FreeSans 6507 0 0 0 io_in_3v3[17]
flabel metal3 s -400 168139 240 168195 0 FreeSans 6507 0 0 0 io_in_3v3[18]
flabel metal3 s -400 146528 240 146584 0 FreeSans 6507 0 0 0 io_in_3v3[19]
flabel metal3 s 291760 3136 292400 3192 0 FreeSans 6507 0 0 0 io_in_3v3[1]
flabel metal3 s -400 125017 240 125073 0 FreeSans 6507 0 0 0 io_in_3v3[20]
flabel metal3 s -400 61206 240 61262 0 FreeSans 6507 0 0 0 io_in_3v3[21]
flabel metal3 s -400 39595 240 39651 0 FreeSans 6507 0 0 0 io_in_3v3[22]
flabel metal3 s -400 17984 240 18040 0 FreeSans 6507 0 0 0 io_in_3v3[23]
flabel metal3 s -400 7273 240 7329 0 FreeSans 6507 0 0 0 io_in_3v3[24]
flabel metal3 s -400 4909 240 4965 0 FreeSans 6507 0 0 0 io_in_3v3[25]
flabel metal3 s -400 2545 240 2601 0 FreeSans 6507 0 0 0 io_in_3v3[26]
flabel metal3 s 291760 5500 292400 5556 0 FreeSans 6507 0 0 0 io_in_3v3[2]
flabel metal3 s 291760 7864 292400 7920 0 FreeSans 6507 0 0 0 io_in_3v3[3]
flabel metal3 s 291760 10228 292400 10284 0 FreeSans 6507 0 0 0 io_in_3v3[4]
flabel metal3 s 291760 23457 292400 23513 0 FreeSans 6507 0 0 0 io_in_3v3[5]
flabel metal3 s 291760 45786 292400 45842 0 FreeSans 6507 0 0 0 io_in_3v3[6]
flabel metal3 s 291760 135797 292400 135853 0 FreeSans 6507 0 0 0 io_in_3v3[7]
flabel metal3 s 291760 158008 292400 158064 0 FreeSans 6507 0 0 0 io_in_3v3[8]
flabel metal3 s 291760 180619 292400 180675 0 FreeSans 6507 0 0 0 io_in_3v3[9]
flabel metal3 s 291760 2545 292400 2601 0 FreeSans 6507 0 0 0 io_oeb[0]
flabel metal3 s 291760 205603 292400 205659 0 FreeSans 6507 0 0 0 io_oeb[10]
flabel metal3 s 291760 227814 292400 227870 0 FreeSans 6507 0 0 0 io_oeb[11]
flabel metal3 s 291760 250025 292400 250081 0 FreeSans 6507 0 0 0 io_oeb[12]
flabel metal3 s 291760 294736 292400 294792 0 FreeSans 6507 0 0 0 io_oeb[13]
flabel metal3 s -400 252810 240 252866 0 FreeSans 6507 0 0 0 io_oeb[14]
flabel metal3 s -400 231199 240 231255 0 FreeSans 6507 0 0 0 io_oeb[15]
flabel metal3 s -400 209588 240 209644 0 FreeSans 6507 0 0 0 io_oeb[16]
flabel metal3 s -400 187977 240 188033 0 FreeSans 6507 0 0 0 io_oeb[17]
flabel metal3 s -400 166366 240 166422 0 FreeSans 6507 0 0 0 io_oeb[18]
flabel metal3 s -400 144755 240 144811 0 FreeSans 6507 0 0 0 io_oeb[19]
flabel metal3 s 291760 4909 292400 4965 0 FreeSans 6507 0 0 0 io_oeb[1]
flabel metal3 s -400 123244 240 123300 0 FreeSans 6507 0 0 0 io_oeb[20]
flabel metal3 s -400 59433 240 59489 0 FreeSans 6507 0 0 0 io_oeb[21]
flabel metal3 s -400 37822 240 37878 0 FreeSans 6507 0 0 0 io_oeb[22]
flabel metal3 s -400 16211 240 16267 0 FreeSans 6507 0 0 0 io_oeb[23]
flabel metal3 s -400 5500 240 5556 0 FreeSans 6507 0 0 0 io_oeb[24]
flabel metal3 s -400 3136 240 3192 0 FreeSans 6507 0 0 0 io_oeb[25]
flabel metal3 s -400 772 240 828 0 FreeSans 6507 0 0 0 io_oeb[26]
flabel metal3 s 291760 7273 292400 7329 0 FreeSans 6507 0 0 0 io_oeb[2]
flabel metal3 s 291760 9637 292400 9693 0 FreeSans 6507 0 0 0 io_oeb[3]
flabel metal3 s 291760 12001 292400 12057 0 FreeSans 6507 0 0 0 io_oeb[4]
flabel metal3 s 291760 25230 292400 25286 0 FreeSans 6507 0 0 0 io_oeb[5]
flabel metal3 s 291760 47559 292400 47615 0 FreeSans 6507 0 0 0 io_oeb[6]
flabel metal3 s 291760 137570 292400 137626 0 FreeSans 6507 0 0 0 io_oeb[7]
flabel metal3 s 291760 159781 292400 159837 0 FreeSans 6507 0 0 0 io_oeb[8]
flabel metal3 s 291760 182392 292400 182448 0 FreeSans 6507 0 0 0 io_oeb[9]
flabel metal3 s 291760 1954 292400 2010 0 FreeSans 6507 0 0 0 io_out[0]
flabel metal3 s 291760 205012 292400 205068 0 FreeSans 6507 0 0 0 io_out[10]
flabel metal3 s 291760 227223 292400 227279 0 FreeSans 6507 0 0 0 io_out[11]
flabel metal3 s 291760 249434 292400 249490 0 FreeSans 6507 0 0 0 io_out[12]
flabel metal3 s 291760 294145 292400 294201 0 FreeSans 6507 0 0 0 io_out[13]
flabel metal3 s -400 253401 240 253457 0 FreeSans 6507 0 0 0 io_out[14]
flabel metal3 s -400 231790 240 231846 0 FreeSans 6507 0 0 0 io_out[15]
flabel metal3 s -400 210179 240 210235 0 FreeSans 6507 0 0 0 io_out[16]
flabel metal3 s -400 188568 240 188624 0 FreeSans 6507 0 0 0 io_out[17]
flabel metal3 s -400 166957 240 167013 0 FreeSans 6507 0 0 0 io_out[18]
flabel metal3 s -400 145346 240 145402 0 FreeSans 6507 0 0 0 io_out[19]
flabel metal3 s 291760 4318 292400 4374 0 FreeSans 6507 0 0 0 io_out[1]
flabel metal3 s -400 123835 240 123891 0 FreeSans 6507 0 0 0 io_out[20]
flabel metal3 s -400 60024 240 60080 0 FreeSans 6507 0 0 0 io_out[21]
flabel metal3 s -400 38413 240 38469 0 FreeSans 6507 0 0 0 io_out[22]
flabel metal3 s -400 16802 240 16858 0 FreeSans 6507 0 0 0 io_out[23]
flabel metal3 s -400 6091 240 6147 0 FreeSans 6507 0 0 0 io_out[24]
flabel metal3 s -400 3727 240 3783 0 FreeSans 6507 0 0 0 io_out[25]
flabel metal3 s -400 1363 240 1419 0 FreeSans 6507 0 0 0 io_out[26]
flabel metal3 s 291760 6682 292400 6738 0 FreeSans 6507 0 0 0 io_out[2]
flabel metal3 s 291760 9046 292400 9102 0 FreeSans 6507 0 0 0 io_out[3]
flabel metal3 s 291760 11410 292400 11466 0 FreeSans 6507 0 0 0 io_out[4]
flabel metal3 s 291760 24639 292400 24695 0 FreeSans 6507 0 0 0 io_out[5]
flabel metal3 s 291760 46968 292400 47024 0 FreeSans 6507 0 0 0 io_out[6]
flabel metal3 s 291760 136979 292400 137035 0 FreeSans 6507 0 0 0 io_out[7]
flabel metal3 s 291760 159190 292400 159246 0 FreeSans 6507 0 0 0 io_out[8]
flabel metal3 s 291760 181801 292400 181857 0 FreeSans 6507 0 0 0 io_out[9]
flabel metal2 s 62908 -400 62964 240 0 FreeSans 6507 90 0 0 la_data_in[0]
flabel metal2 s 240208 -400 240264 240 0 FreeSans 6507 90 0 0 la_data_in[100]
flabel metal2 s 241981 -400 242037 240 0 FreeSans 6507 90 0 0 la_data_in[101]
flabel metal2 s 243754 -400 243810 240 0 FreeSans 6507 90 0 0 la_data_in[102]
flabel metal2 s 245527 -400 245583 240 0 FreeSans 6507 90 0 0 la_data_in[103]
flabel metal2 s 247300 -400 247356 240 0 FreeSans 6507 90 0 0 la_data_in[104]
flabel metal2 s 249073 -400 249129 240 0 FreeSans 6507 90 0 0 la_data_in[105]
flabel metal2 s 250846 -400 250902 240 0 FreeSans 6507 90 0 0 la_data_in[106]
flabel metal2 s 252619 -400 252675 240 0 FreeSans 6507 90 0 0 la_data_in[107]
flabel metal2 s 254392 -400 254448 240 0 FreeSans 6507 90 0 0 la_data_in[108]
flabel metal2 s 256165 -400 256221 240 0 FreeSans 6507 90 0 0 la_data_in[109]
flabel metal2 s 80638 -400 80694 240 0 FreeSans 6507 90 0 0 la_data_in[10]
flabel metal2 s 257938 -400 257994 240 0 FreeSans 6507 90 0 0 la_data_in[110]
flabel metal2 s 259711 -400 259767 240 0 FreeSans 6507 90 0 0 la_data_in[111]
flabel metal2 s 261484 -400 261540 240 0 FreeSans 6507 90 0 0 la_data_in[112]
flabel metal2 s 263257 -400 263313 240 0 FreeSans 6507 90 0 0 la_data_in[113]
flabel metal2 s 265030 -400 265086 240 0 FreeSans 6507 90 0 0 la_data_in[114]
flabel metal2 s 266803 -400 266859 240 0 FreeSans 6507 90 0 0 la_data_in[115]
flabel metal2 s 268576 -400 268632 240 0 FreeSans 6507 90 0 0 la_data_in[116]
flabel metal2 s 270349 -400 270405 240 0 FreeSans 6507 90 0 0 la_data_in[117]
flabel metal2 s 272122 -400 272178 240 0 FreeSans 6507 90 0 0 la_data_in[118]
flabel metal2 s 273895 -400 273951 240 0 FreeSans 6507 90 0 0 la_data_in[119]
flabel metal2 s 82411 -400 82467 240 0 FreeSans 6507 90 0 0 la_data_in[11]
flabel metal2 s 275668 -400 275724 240 0 FreeSans 6507 90 0 0 la_data_in[120]
flabel metal2 s 277441 -400 277497 240 0 FreeSans 6507 90 0 0 la_data_in[121]
flabel metal2 s 279214 -400 279270 240 0 FreeSans 6507 90 0 0 la_data_in[122]
flabel metal2 s 280987 -400 281043 240 0 FreeSans 6507 90 0 0 la_data_in[123]
flabel metal2 s 282760 -400 282816 240 0 FreeSans 6507 90 0 0 la_data_in[124]
flabel metal2 s 284533 -400 284589 240 0 FreeSans 6507 90 0 0 la_data_in[125]
flabel metal2 s 286306 -400 286362 240 0 FreeSans 6507 90 0 0 la_data_in[126]
flabel metal2 s 288079 -400 288135 240 0 FreeSans 6507 90 0 0 la_data_in[127]
flabel metal2 s 84184 -400 84240 240 0 FreeSans 6507 90 0 0 la_data_in[12]
flabel metal2 s 85957 -400 86013 240 0 FreeSans 6507 90 0 0 la_data_in[13]
flabel metal2 s 87730 -400 87786 240 0 FreeSans 6507 90 0 0 la_data_in[14]
flabel metal2 s 89503 -400 89559 240 0 FreeSans 6507 90 0 0 la_data_in[15]
flabel metal2 s 91276 -400 91332 240 0 FreeSans 6507 90 0 0 la_data_in[16]
flabel metal2 s 93049 -400 93105 240 0 FreeSans 6507 90 0 0 la_data_in[17]
flabel metal2 s 94822 -400 94878 240 0 FreeSans 6507 90 0 0 la_data_in[18]
flabel metal2 s 96595 -400 96651 240 0 FreeSans 6507 90 0 0 la_data_in[19]
flabel metal2 s 64681 -400 64737 240 0 FreeSans 6507 90 0 0 la_data_in[1]
flabel metal2 s 98368 -400 98424 240 0 FreeSans 6507 90 0 0 la_data_in[20]
flabel metal2 s 100141 -400 100197 240 0 FreeSans 6507 90 0 0 la_data_in[21]
flabel metal2 s 101914 -400 101970 240 0 FreeSans 6507 90 0 0 la_data_in[22]
flabel metal2 s 103687 -400 103743 240 0 FreeSans 6507 90 0 0 la_data_in[23]
flabel metal2 s 105460 -400 105516 240 0 FreeSans 6507 90 0 0 la_data_in[24]
flabel metal2 s 107233 -400 107289 240 0 FreeSans 6507 90 0 0 la_data_in[25]
flabel metal2 s 109006 -400 109062 240 0 FreeSans 6507 90 0 0 la_data_in[26]
flabel metal2 s 110779 -400 110835 240 0 FreeSans 6507 90 0 0 la_data_in[27]
flabel metal2 s 112552 -400 112608 240 0 FreeSans 6507 90 0 0 la_data_in[28]
flabel metal2 s 114325 -400 114381 240 0 FreeSans 6507 90 0 0 la_data_in[29]
flabel metal2 s 66454 -400 66510 240 0 FreeSans 6507 90 0 0 la_data_in[2]
flabel metal2 s 116098 -400 116154 240 0 FreeSans 6507 90 0 0 la_data_in[30]
flabel metal2 s 117871 -400 117927 240 0 FreeSans 6507 90 0 0 la_data_in[31]
flabel metal2 s 119644 -400 119700 240 0 FreeSans 6507 90 0 0 la_data_in[32]
flabel metal2 s 121417 -400 121473 240 0 FreeSans 6507 90 0 0 la_data_in[33]
flabel metal2 s 123190 -400 123246 240 0 FreeSans 6507 90 0 0 la_data_in[34]
flabel metal2 s 124963 -400 125019 240 0 FreeSans 6507 90 0 0 la_data_in[35]
flabel metal2 s 126736 -400 126792 240 0 FreeSans 6507 90 0 0 la_data_in[36]
flabel metal2 s 128509 -400 128565 240 0 FreeSans 6507 90 0 0 la_data_in[37]
flabel metal2 s 130282 -400 130338 240 0 FreeSans 6507 90 0 0 la_data_in[38]
flabel metal2 s 132055 -400 132111 240 0 FreeSans 6507 90 0 0 la_data_in[39]
flabel metal2 s 68227 -400 68283 240 0 FreeSans 6507 90 0 0 la_data_in[3]
flabel metal2 s 133828 -400 133884 240 0 FreeSans 6507 90 0 0 la_data_in[40]
flabel metal2 s 135601 -400 135657 240 0 FreeSans 6507 90 0 0 la_data_in[41]
flabel metal2 s 137374 -400 137430 240 0 FreeSans 6507 90 0 0 la_data_in[42]
flabel metal2 s 139147 -400 139203 240 0 FreeSans 6507 90 0 0 la_data_in[43]
flabel metal2 s 140920 -400 140976 240 0 FreeSans 6507 90 0 0 la_data_in[44]
flabel metal2 s 142693 -400 142749 240 0 FreeSans 6507 90 0 0 la_data_in[45]
flabel metal2 s 144466 -400 144522 240 0 FreeSans 6507 90 0 0 la_data_in[46]
flabel metal2 s 146239 -400 146295 240 0 FreeSans 6507 90 0 0 la_data_in[47]
flabel metal2 s 148012 -400 148068 240 0 FreeSans 6507 90 0 0 la_data_in[48]
flabel metal2 s 149785 -400 149841 240 0 FreeSans 6507 90 0 0 la_data_in[49]
flabel metal2 s 70000 -400 70056 240 0 FreeSans 6507 90 0 0 la_data_in[4]
flabel metal2 s 151558 -400 151614 240 0 FreeSans 6507 90 0 0 la_data_in[50]
flabel metal2 s 153331 -400 153387 240 0 FreeSans 6507 90 0 0 la_data_in[51]
flabel metal2 s 155104 -400 155160 240 0 FreeSans 6507 90 0 0 la_data_in[52]
flabel metal2 s 156877 -400 156933 240 0 FreeSans 6507 90 0 0 la_data_in[53]
flabel metal2 s 158650 -400 158706 240 0 FreeSans 6507 90 0 0 la_data_in[54]
flabel metal2 s 160423 -400 160479 240 0 FreeSans 6507 90 0 0 la_data_in[55]
flabel metal2 s 162196 -400 162252 240 0 FreeSans 6507 90 0 0 la_data_in[56]
flabel metal2 s 163969 -400 164025 240 0 FreeSans 6507 90 0 0 la_data_in[57]
flabel metal2 s 165742 -400 165798 240 0 FreeSans 6507 90 0 0 la_data_in[58]
flabel metal2 s 167515 -400 167571 240 0 FreeSans 6507 90 0 0 la_data_in[59]
flabel metal2 s 71773 -400 71829 240 0 FreeSans 6507 90 0 0 la_data_in[5]
flabel metal2 s 169288 -400 169344 240 0 FreeSans 6507 90 0 0 la_data_in[60]
flabel metal2 s 171061 -400 171117 240 0 FreeSans 6507 90 0 0 la_data_in[61]
flabel metal2 s 172834 -400 172890 240 0 FreeSans 6507 90 0 0 la_data_in[62]
flabel metal2 s 174607 -400 174663 240 0 FreeSans 6507 90 0 0 la_data_in[63]
flabel metal2 s 176380 -400 176436 240 0 FreeSans 6507 90 0 0 la_data_in[64]
flabel metal2 s 178153 -400 178209 240 0 FreeSans 6507 90 0 0 la_data_in[65]
flabel metal2 s 179926 -400 179982 240 0 FreeSans 6507 90 0 0 la_data_in[66]
flabel metal2 s 181699 -400 181755 240 0 FreeSans 6507 90 0 0 la_data_in[67]
flabel metal2 s 183472 -400 183528 240 0 FreeSans 6507 90 0 0 la_data_in[68]
flabel metal2 s 185245 -400 185301 240 0 FreeSans 6507 90 0 0 la_data_in[69]
flabel metal2 s 73546 -400 73602 240 0 FreeSans 6507 90 0 0 la_data_in[6]
flabel metal2 s 187018 -400 187074 240 0 FreeSans 6507 90 0 0 la_data_in[70]
flabel metal2 s 188791 -400 188847 240 0 FreeSans 6507 90 0 0 la_data_in[71]
flabel metal2 s 190564 -400 190620 240 0 FreeSans 6507 90 0 0 la_data_in[72]
flabel metal2 s 192337 -400 192393 240 0 FreeSans 6507 90 0 0 la_data_in[73]
flabel metal2 s 194110 -400 194166 240 0 FreeSans 6507 90 0 0 la_data_in[74]
flabel metal2 s 195883 -400 195939 240 0 FreeSans 6507 90 0 0 la_data_in[75]
flabel metal2 s 197656 -400 197712 240 0 FreeSans 6507 90 0 0 la_data_in[76]
flabel metal2 s 199429 -400 199485 240 0 FreeSans 6507 90 0 0 la_data_in[77]
flabel metal2 s 201202 -400 201258 240 0 FreeSans 6507 90 0 0 la_data_in[78]
flabel metal2 s 202975 -400 203031 240 0 FreeSans 6507 90 0 0 la_data_in[79]
flabel metal2 s 75319 -400 75375 240 0 FreeSans 6507 90 0 0 la_data_in[7]
flabel metal2 s 204748 -400 204804 240 0 FreeSans 6507 90 0 0 la_data_in[80]
flabel metal2 s 206521 -400 206577 240 0 FreeSans 6507 90 0 0 la_data_in[81]
flabel metal2 s 208294 -400 208350 240 0 FreeSans 6507 90 0 0 la_data_in[82]
flabel metal2 s 210067 -400 210123 240 0 FreeSans 6507 90 0 0 la_data_in[83]
flabel metal2 s 211840 -400 211896 240 0 FreeSans 6507 90 0 0 la_data_in[84]
flabel metal2 s 213613 -400 213669 240 0 FreeSans 6507 90 0 0 la_data_in[85]
flabel metal2 s 215386 -400 215442 240 0 FreeSans 6507 90 0 0 la_data_in[86]
flabel metal2 s 217159 -400 217215 240 0 FreeSans 6507 90 0 0 la_data_in[87]
flabel metal2 s 218932 -400 218988 240 0 FreeSans 6507 90 0 0 la_data_in[88]
flabel metal2 s 220705 -400 220761 240 0 FreeSans 6507 90 0 0 la_data_in[89]
flabel metal2 s 77092 -400 77148 240 0 FreeSans 6507 90 0 0 la_data_in[8]
flabel metal2 s 222478 -400 222534 240 0 FreeSans 6507 90 0 0 la_data_in[90]
flabel metal2 s 224251 -400 224307 240 0 FreeSans 6507 90 0 0 la_data_in[91]
flabel metal2 s 226024 -400 226080 240 0 FreeSans 6507 90 0 0 la_data_in[92]
flabel metal2 s 227797 -400 227853 240 0 FreeSans 6507 90 0 0 la_data_in[93]
flabel metal2 s 229570 -400 229626 240 0 FreeSans 6507 90 0 0 la_data_in[94]
flabel metal2 s 231343 -400 231399 240 0 FreeSans 6507 90 0 0 la_data_in[95]
flabel metal2 s 233116 -400 233172 240 0 FreeSans 6507 90 0 0 la_data_in[96]
flabel metal2 s 234889 -400 234945 240 0 FreeSans 6507 90 0 0 la_data_in[97]
flabel metal2 s 236662 -400 236718 240 0 FreeSans 6507 90 0 0 la_data_in[98]
flabel metal2 s 238435 -400 238491 240 0 FreeSans 6507 90 0 0 la_data_in[99]
flabel metal2 s 78865 -400 78921 240 0 FreeSans 6507 90 0 0 la_data_in[9]
flabel metal2 s 63499 -400 63555 240 0 FreeSans 6507 90 0 0 la_data_out[0]
flabel metal2 s 240799 -400 240855 240 0 FreeSans 6507 90 0 0 la_data_out[100]
flabel metal2 s 242572 -400 242628 240 0 FreeSans 6507 90 0 0 la_data_out[101]
flabel metal2 s 244345 -400 244401 240 0 FreeSans 6507 90 0 0 la_data_out[102]
flabel metal2 s 246118 -400 246174 240 0 FreeSans 6507 90 0 0 la_data_out[103]
flabel metal2 s 247891 -400 247947 240 0 FreeSans 6507 90 0 0 la_data_out[104]
flabel metal2 s 249664 -400 249720 240 0 FreeSans 6507 90 0 0 la_data_out[105]
flabel metal2 s 251437 -400 251493 240 0 FreeSans 6507 90 0 0 la_data_out[106]
flabel metal2 s 253210 -400 253266 240 0 FreeSans 6507 90 0 0 la_data_out[107]
flabel metal2 s 254983 -400 255039 240 0 FreeSans 6507 90 0 0 la_data_out[108]
flabel metal2 s 256756 -400 256812 240 0 FreeSans 6507 90 0 0 la_data_out[109]
flabel metal2 s 81229 -400 81285 240 0 FreeSans 6507 90 0 0 la_data_out[10]
flabel metal2 s 258529 -400 258585 240 0 FreeSans 6507 90 0 0 la_data_out[110]
flabel metal2 s 260302 -400 260358 240 0 FreeSans 6507 90 0 0 la_data_out[111]
flabel metal2 s 262075 -400 262131 240 0 FreeSans 6507 90 0 0 la_data_out[112]
flabel metal2 s 263848 -400 263904 240 0 FreeSans 6507 90 0 0 la_data_out[113]
flabel metal2 s 265621 -400 265677 240 0 FreeSans 6507 90 0 0 la_data_out[114]
flabel metal2 s 267394 -400 267450 240 0 FreeSans 6507 90 0 0 la_data_out[115]
flabel metal2 s 269167 -400 269223 240 0 FreeSans 6507 90 0 0 la_data_out[116]
flabel metal2 s 270940 -400 270996 240 0 FreeSans 6507 90 0 0 la_data_out[117]
flabel metal2 s 272713 -400 272769 240 0 FreeSans 6507 90 0 0 la_data_out[118]
flabel metal2 s 274486 -400 274542 240 0 FreeSans 6507 90 0 0 la_data_out[119]
flabel metal2 s 83002 -400 83058 240 0 FreeSans 6507 90 0 0 la_data_out[11]
flabel metal2 s 276259 -400 276315 240 0 FreeSans 6507 90 0 0 la_data_out[120]
flabel metal2 s 278032 -400 278088 240 0 FreeSans 6507 90 0 0 la_data_out[121]
flabel metal2 s 279805 -400 279861 240 0 FreeSans 6507 90 0 0 la_data_out[122]
flabel metal2 s 281578 -400 281634 240 0 FreeSans 6507 90 0 0 la_data_out[123]
flabel metal2 s 283351 -400 283407 240 0 FreeSans 6507 90 0 0 la_data_out[124]
flabel metal2 s 285124 -400 285180 240 0 FreeSans 6507 90 0 0 la_data_out[125]
flabel metal2 s 286897 -400 286953 240 0 FreeSans 6507 90 0 0 la_data_out[126]
flabel metal2 s 288670 -400 288726 240 0 FreeSans 6507 90 0 0 la_data_out[127]
flabel metal2 s 84775 -400 84831 240 0 FreeSans 6507 90 0 0 la_data_out[12]
flabel metal2 s 86548 -400 86604 240 0 FreeSans 6507 90 0 0 la_data_out[13]
flabel metal2 s 88321 -400 88377 240 0 FreeSans 6507 90 0 0 la_data_out[14]
flabel metal2 s 90094 -400 90150 240 0 FreeSans 6507 90 0 0 la_data_out[15]
flabel metal2 s 91867 -400 91923 240 0 FreeSans 6507 90 0 0 la_data_out[16]
flabel metal2 s 93640 -400 93696 240 0 FreeSans 6507 90 0 0 la_data_out[17]
flabel metal2 s 95413 -400 95469 240 0 FreeSans 6507 90 0 0 la_data_out[18]
flabel metal2 s 97186 -400 97242 240 0 FreeSans 6507 90 0 0 la_data_out[19]
flabel metal2 s 65272 -400 65328 240 0 FreeSans 6507 90 0 0 la_data_out[1]
flabel metal2 s 98959 -400 99015 240 0 FreeSans 6507 90 0 0 la_data_out[20]
flabel metal2 s 100732 -400 100788 240 0 FreeSans 6507 90 0 0 la_data_out[21]
flabel metal2 s 102505 -400 102561 240 0 FreeSans 6507 90 0 0 la_data_out[22]
flabel metal2 s 104278 -400 104334 240 0 FreeSans 6507 90 0 0 la_data_out[23]
flabel metal2 s 106051 -400 106107 240 0 FreeSans 6507 90 0 0 la_data_out[24]
flabel metal2 s 107824 -400 107880 240 0 FreeSans 6507 90 0 0 la_data_out[25]
flabel metal2 s 109597 -400 109653 240 0 FreeSans 6507 90 0 0 la_data_out[26]
flabel metal2 s 111370 -400 111426 240 0 FreeSans 6507 90 0 0 la_data_out[27]
flabel metal2 s 113143 -400 113199 240 0 FreeSans 6507 90 0 0 la_data_out[28]
flabel metal2 s 114916 -400 114972 240 0 FreeSans 6507 90 0 0 la_data_out[29]
flabel metal2 s 67045 -400 67101 240 0 FreeSans 6507 90 0 0 la_data_out[2]
flabel metal2 s 116689 -400 116745 240 0 FreeSans 6507 90 0 0 la_data_out[30]
flabel metal2 s 118462 -400 118518 240 0 FreeSans 6507 90 0 0 la_data_out[31]
flabel metal2 s 120235 -400 120291 240 0 FreeSans 6507 90 0 0 la_data_out[32]
flabel metal2 s 122008 -400 122064 240 0 FreeSans 6507 90 0 0 la_data_out[33]
flabel metal2 s 123781 -400 123837 240 0 FreeSans 6507 90 0 0 la_data_out[34]
flabel metal2 s 125554 -400 125610 240 0 FreeSans 6507 90 0 0 la_data_out[35]
flabel metal2 s 127327 -400 127383 240 0 FreeSans 6507 90 0 0 la_data_out[36]
flabel metal2 s 129100 -400 129156 240 0 FreeSans 6507 90 0 0 la_data_out[37]
flabel metal2 s 130873 -400 130929 240 0 FreeSans 6507 90 0 0 la_data_out[38]
flabel metal2 s 132646 -400 132702 240 0 FreeSans 6507 90 0 0 la_data_out[39]
flabel metal2 s 68818 -400 68874 240 0 FreeSans 6507 90 0 0 la_data_out[3]
flabel metal2 s 134419 -400 134475 240 0 FreeSans 6507 90 0 0 la_data_out[40]
flabel metal2 s 136192 -400 136248 240 0 FreeSans 6507 90 0 0 la_data_out[41]
flabel metal2 s 137965 -400 138021 240 0 FreeSans 6507 90 0 0 la_data_out[42]
flabel metal2 s 139738 -400 139794 240 0 FreeSans 6507 90 0 0 la_data_out[43]
flabel metal2 s 141511 -400 141567 240 0 FreeSans 6507 90 0 0 la_data_out[44]
flabel metal2 s 143284 -400 143340 240 0 FreeSans 6507 90 0 0 la_data_out[45]
flabel metal2 s 145057 -400 145113 240 0 FreeSans 6507 90 0 0 la_data_out[46]
flabel metal2 s 146830 -400 146886 240 0 FreeSans 6507 90 0 0 la_data_out[47]
flabel metal2 s 148603 -400 148659 240 0 FreeSans 6507 90 0 0 la_data_out[48]
flabel metal2 s 150376 -400 150432 240 0 FreeSans 6507 90 0 0 la_data_out[49]
flabel metal2 s 70591 -400 70647 240 0 FreeSans 6507 90 0 0 la_data_out[4]
flabel metal2 s 152149 -400 152205 240 0 FreeSans 6507 90 0 0 la_data_out[50]
flabel metal2 s 153922 -400 153978 240 0 FreeSans 6507 90 0 0 la_data_out[51]
flabel metal2 s 155695 -400 155751 240 0 FreeSans 6507 90 0 0 la_data_out[52]
flabel metal2 s 157468 -400 157524 240 0 FreeSans 6507 90 0 0 la_data_out[53]
flabel metal2 s 159241 -400 159297 240 0 FreeSans 6507 90 0 0 la_data_out[54]
flabel metal2 s 161014 -400 161070 240 0 FreeSans 6507 90 0 0 la_data_out[55]
flabel metal2 s 162787 -400 162843 240 0 FreeSans 6507 90 0 0 la_data_out[56]
flabel metal2 s 164560 -400 164616 240 0 FreeSans 6507 90 0 0 la_data_out[57]
flabel metal2 s 166333 -400 166389 240 0 FreeSans 6507 90 0 0 la_data_out[58]
flabel metal2 s 168106 -400 168162 240 0 FreeSans 6507 90 0 0 la_data_out[59]
flabel metal2 s 72364 -400 72420 240 0 FreeSans 6507 90 0 0 la_data_out[5]
flabel metal2 s 169879 -400 169935 240 0 FreeSans 6507 90 0 0 la_data_out[60]
flabel metal2 s 171652 -400 171708 240 0 FreeSans 6507 90 0 0 la_data_out[61]
flabel metal2 s 173425 -400 173481 240 0 FreeSans 6507 90 0 0 la_data_out[62]
flabel metal2 s 175198 -400 175254 240 0 FreeSans 6507 90 0 0 la_data_out[63]
flabel metal2 s 176971 -400 177027 240 0 FreeSans 6507 90 0 0 la_data_out[64]
flabel metal2 s 178744 -400 178800 240 0 FreeSans 6507 90 0 0 la_data_out[65]
flabel metal2 s 180517 -400 180573 240 0 FreeSans 6507 90 0 0 la_data_out[66]
flabel metal2 s 182290 -400 182346 240 0 FreeSans 6507 90 0 0 la_data_out[67]
flabel metal2 s 184063 -400 184119 240 0 FreeSans 6507 90 0 0 la_data_out[68]
flabel metal2 s 185836 -400 185892 240 0 FreeSans 6507 90 0 0 la_data_out[69]
flabel metal2 s 74137 -400 74193 240 0 FreeSans 6507 90 0 0 la_data_out[6]
flabel metal2 s 187609 -400 187665 240 0 FreeSans 6507 90 0 0 la_data_out[70]
flabel metal2 s 189382 -400 189438 240 0 FreeSans 6507 90 0 0 la_data_out[71]
flabel metal2 s 191155 -400 191211 240 0 FreeSans 6507 90 0 0 la_data_out[72]
flabel metal2 s 192928 -400 192984 240 0 FreeSans 6507 90 0 0 la_data_out[73]
flabel metal2 s 194701 -400 194757 240 0 FreeSans 6507 90 0 0 la_data_out[74]
flabel metal2 s 196474 -400 196530 240 0 FreeSans 6507 90 0 0 la_data_out[75]
flabel metal2 s 198247 -400 198303 240 0 FreeSans 6507 90 0 0 la_data_out[76]
flabel metal2 s 200020 -400 200076 240 0 FreeSans 6507 90 0 0 la_data_out[77]
flabel metal2 s 201793 -400 201849 240 0 FreeSans 6507 90 0 0 la_data_out[78]
flabel metal2 s 203566 -400 203622 240 0 FreeSans 6507 90 0 0 la_data_out[79]
flabel metal2 s 75910 -400 75966 240 0 FreeSans 6507 90 0 0 la_data_out[7]
flabel metal2 s 205339 -400 205395 240 0 FreeSans 6507 90 0 0 la_data_out[80]
flabel metal2 s 207112 -400 207168 240 0 FreeSans 6507 90 0 0 la_data_out[81]
flabel metal2 s 208885 -400 208941 240 0 FreeSans 6507 90 0 0 la_data_out[82]
flabel metal2 s 210658 -400 210714 240 0 FreeSans 6507 90 0 0 la_data_out[83]
flabel metal2 s 212431 -400 212487 240 0 FreeSans 6507 90 0 0 la_data_out[84]
flabel metal2 s 214204 -400 214260 240 0 FreeSans 6507 90 0 0 la_data_out[85]
flabel metal2 s 215977 -400 216033 240 0 FreeSans 6507 90 0 0 la_data_out[86]
flabel metal2 s 217750 -400 217806 240 0 FreeSans 6507 90 0 0 la_data_out[87]
flabel metal2 s 219523 -400 219579 240 0 FreeSans 6507 90 0 0 la_data_out[88]
flabel metal2 s 221296 -400 221352 240 0 FreeSans 6507 90 0 0 la_data_out[89]
flabel metal2 s 77683 -400 77739 240 0 FreeSans 6507 90 0 0 la_data_out[8]
flabel metal2 s 223069 -400 223125 240 0 FreeSans 6507 90 0 0 la_data_out[90]
flabel metal2 s 224842 -400 224898 240 0 FreeSans 6507 90 0 0 la_data_out[91]
flabel metal2 s 226615 -400 226671 240 0 FreeSans 6507 90 0 0 la_data_out[92]
flabel metal2 s 228388 -400 228444 240 0 FreeSans 6507 90 0 0 la_data_out[93]
flabel metal2 s 230161 -400 230217 240 0 FreeSans 6507 90 0 0 la_data_out[94]
flabel metal2 s 231934 -400 231990 240 0 FreeSans 6507 90 0 0 la_data_out[95]
flabel metal2 s 233707 -400 233763 240 0 FreeSans 6507 90 0 0 la_data_out[96]
flabel metal2 s 235480 -400 235536 240 0 FreeSans 6507 90 0 0 la_data_out[97]
flabel metal2 s 237253 -400 237309 240 0 FreeSans 6507 90 0 0 la_data_out[98]
flabel metal2 s 239026 -400 239082 240 0 FreeSans 6507 90 0 0 la_data_out[99]
flabel metal2 s 79456 -400 79512 240 0 FreeSans 6507 90 0 0 la_data_out[9]
flabel metal2 s 64090 -400 64146 240 0 FreeSans 6507 90 0 0 la_oenb[0]
flabel metal2 s 241390 -400 241446 240 0 FreeSans 6507 90 0 0 la_oenb[100]
flabel metal2 s 243163 -400 243219 240 0 FreeSans 6507 90 0 0 la_oenb[101]
flabel metal2 s 244936 -400 244992 240 0 FreeSans 6507 90 0 0 la_oenb[102]
flabel metal2 s 246709 -400 246765 240 0 FreeSans 6507 90 0 0 la_oenb[103]
flabel metal2 s 248482 -400 248538 240 0 FreeSans 6507 90 0 0 la_oenb[104]
flabel metal2 s 250255 -400 250311 240 0 FreeSans 6507 90 0 0 la_oenb[105]
flabel metal2 s 252028 -400 252084 240 0 FreeSans 6507 90 0 0 la_oenb[106]
flabel metal2 s 253801 -400 253857 240 0 FreeSans 6507 90 0 0 la_oenb[107]
flabel metal2 s 255574 -400 255630 240 0 FreeSans 6507 90 0 0 la_oenb[108]
flabel metal2 s 257347 -400 257403 240 0 FreeSans 6507 90 0 0 la_oenb[109]
flabel metal2 s 81820 -400 81876 240 0 FreeSans 6507 90 0 0 la_oenb[10]
flabel metal2 s 259120 -400 259176 240 0 FreeSans 6507 90 0 0 la_oenb[110]
flabel metal2 s 260893 -400 260949 240 0 FreeSans 6507 90 0 0 la_oenb[111]
flabel metal2 s 262666 -400 262722 240 0 FreeSans 6507 90 0 0 la_oenb[112]
flabel metal2 s 264439 -400 264495 240 0 FreeSans 6507 90 0 0 la_oenb[113]
flabel metal2 s 266212 -400 266268 240 0 FreeSans 6507 90 0 0 la_oenb[114]
flabel metal2 s 267985 -400 268041 240 0 FreeSans 6507 90 0 0 la_oenb[115]
flabel metal2 s 269758 -400 269814 240 0 FreeSans 6507 90 0 0 la_oenb[116]
flabel metal2 s 271531 -400 271587 240 0 FreeSans 6507 90 0 0 la_oenb[117]
flabel metal2 s 273304 -400 273360 240 0 FreeSans 6507 90 0 0 la_oenb[118]
flabel metal2 s 275077 -400 275133 240 0 FreeSans 6507 90 0 0 la_oenb[119]
flabel metal2 s 83593 -400 83649 240 0 FreeSans 6507 90 0 0 la_oenb[11]
flabel metal2 s 276850 -400 276906 240 0 FreeSans 6507 90 0 0 la_oenb[120]
flabel metal2 s 278623 -400 278679 240 0 FreeSans 6507 90 0 0 la_oenb[121]
flabel metal2 s 280396 -400 280452 240 0 FreeSans 6507 90 0 0 la_oenb[122]
flabel metal2 s 282169 -400 282225 240 0 FreeSans 6507 90 0 0 la_oenb[123]
flabel metal2 s 283942 -400 283998 240 0 FreeSans 6507 90 0 0 la_oenb[124]
flabel metal2 s 285715 -400 285771 240 0 FreeSans 6507 90 0 0 la_oenb[125]
flabel metal2 s 287488 -400 287544 240 0 FreeSans 6507 90 0 0 la_oenb[126]
flabel metal2 s 289261 -400 289317 240 0 FreeSans 6507 90 0 0 la_oenb[127]
flabel metal2 s 85366 -400 85422 240 0 FreeSans 6507 90 0 0 la_oenb[12]
flabel metal2 s 87139 -400 87195 240 0 FreeSans 6507 90 0 0 la_oenb[13]
flabel metal2 s 88912 -400 88968 240 0 FreeSans 6507 90 0 0 la_oenb[14]
flabel metal2 s 90685 -400 90741 240 0 FreeSans 6507 90 0 0 la_oenb[15]
flabel metal2 s 92458 -400 92514 240 0 FreeSans 6507 90 0 0 la_oenb[16]
flabel metal2 s 94231 -400 94287 240 0 FreeSans 6507 90 0 0 la_oenb[17]
flabel metal2 s 96004 -400 96060 240 0 FreeSans 6507 90 0 0 la_oenb[18]
flabel metal2 s 97777 -400 97833 240 0 FreeSans 6507 90 0 0 la_oenb[19]
flabel metal2 s 65863 -400 65919 240 0 FreeSans 6507 90 0 0 la_oenb[1]
flabel metal2 s 99550 -400 99606 240 0 FreeSans 6507 90 0 0 la_oenb[20]
flabel metal2 s 101323 -400 101379 240 0 FreeSans 6507 90 0 0 la_oenb[21]
flabel metal2 s 103096 -400 103152 240 0 FreeSans 6507 90 0 0 la_oenb[22]
flabel metal2 s 104869 -400 104925 240 0 FreeSans 6507 90 0 0 la_oenb[23]
flabel metal2 s 106642 -400 106698 240 0 FreeSans 6507 90 0 0 la_oenb[24]
flabel metal2 s 108415 -400 108471 240 0 FreeSans 6507 90 0 0 la_oenb[25]
flabel metal2 s 110188 -400 110244 240 0 FreeSans 6507 90 0 0 la_oenb[26]
flabel metal2 s 111961 -400 112017 240 0 FreeSans 6507 90 0 0 la_oenb[27]
flabel metal2 s 113734 -400 113790 240 0 FreeSans 6507 90 0 0 la_oenb[28]
flabel metal2 s 115507 -400 115563 240 0 FreeSans 6507 90 0 0 la_oenb[29]
flabel metal2 s 67636 -400 67692 240 0 FreeSans 6507 90 0 0 la_oenb[2]
flabel metal2 s 117280 -400 117336 240 0 FreeSans 6507 90 0 0 la_oenb[30]
flabel metal2 s 119053 -400 119109 240 0 FreeSans 6507 90 0 0 la_oenb[31]
flabel metal2 s 120826 -400 120882 240 0 FreeSans 6507 90 0 0 la_oenb[32]
flabel metal2 s 122599 -400 122655 240 0 FreeSans 6507 90 0 0 la_oenb[33]
flabel metal2 s 124372 -400 124428 240 0 FreeSans 6507 90 0 0 la_oenb[34]
flabel metal2 s 126145 -400 126201 240 0 FreeSans 6507 90 0 0 la_oenb[35]
flabel metal2 s 127918 -400 127974 240 0 FreeSans 6507 90 0 0 la_oenb[36]
flabel metal2 s 129691 -400 129747 240 0 FreeSans 6507 90 0 0 la_oenb[37]
flabel metal2 s 131464 -400 131520 240 0 FreeSans 6507 90 0 0 la_oenb[38]
flabel metal2 s 133237 -400 133293 240 0 FreeSans 6507 90 0 0 la_oenb[39]
flabel metal2 s 69409 -400 69465 240 0 FreeSans 6507 90 0 0 la_oenb[3]
flabel metal2 s 135010 -400 135066 240 0 FreeSans 6507 90 0 0 la_oenb[40]
flabel metal2 s 136783 -400 136839 240 0 FreeSans 6507 90 0 0 la_oenb[41]
flabel metal2 s 138556 -400 138612 240 0 FreeSans 6507 90 0 0 la_oenb[42]
flabel metal2 s 140329 -400 140385 240 0 FreeSans 6507 90 0 0 la_oenb[43]
flabel metal2 s 142102 -400 142158 240 0 FreeSans 6507 90 0 0 la_oenb[44]
flabel metal2 s 143875 -400 143931 240 0 FreeSans 6507 90 0 0 la_oenb[45]
flabel metal2 s 145648 -400 145704 240 0 FreeSans 6507 90 0 0 la_oenb[46]
flabel metal2 s 147421 -400 147477 240 0 FreeSans 6507 90 0 0 la_oenb[47]
flabel metal2 s 149194 -400 149250 240 0 FreeSans 6507 90 0 0 la_oenb[48]
flabel metal2 s 150967 -400 151023 240 0 FreeSans 6507 90 0 0 la_oenb[49]
flabel metal2 s 71182 -400 71238 240 0 FreeSans 6507 90 0 0 la_oenb[4]
flabel metal2 s 152740 -400 152796 240 0 FreeSans 6507 90 0 0 la_oenb[50]
flabel metal2 s 154513 -400 154569 240 0 FreeSans 6507 90 0 0 la_oenb[51]
flabel metal2 s 156286 -400 156342 240 0 FreeSans 6507 90 0 0 la_oenb[52]
flabel metal2 s 158059 -400 158115 240 0 FreeSans 6507 90 0 0 la_oenb[53]
flabel metal2 s 159832 -400 159888 240 0 FreeSans 6507 90 0 0 la_oenb[54]
flabel metal2 s 161605 -400 161661 240 0 FreeSans 6507 90 0 0 la_oenb[55]
flabel metal2 s 163378 -400 163434 240 0 FreeSans 6507 90 0 0 la_oenb[56]
flabel metal2 s 165151 -400 165207 240 0 FreeSans 6507 90 0 0 la_oenb[57]
flabel metal2 s 166924 -400 166980 240 0 FreeSans 6507 90 0 0 la_oenb[58]
flabel metal2 s 168697 -400 168753 240 0 FreeSans 6507 90 0 0 la_oenb[59]
flabel metal2 s 72955 -400 73011 240 0 FreeSans 6507 90 0 0 la_oenb[5]
flabel metal2 s 170470 -400 170526 240 0 FreeSans 6507 90 0 0 la_oenb[60]
flabel metal2 s 172243 -400 172299 240 0 FreeSans 6507 90 0 0 la_oenb[61]
flabel metal2 s 174016 -400 174072 240 0 FreeSans 6507 90 0 0 la_oenb[62]
flabel metal2 s 175789 -400 175845 240 0 FreeSans 6507 90 0 0 la_oenb[63]
flabel metal2 s 177562 -400 177618 240 0 FreeSans 6507 90 0 0 la_oenb[64]
flabel metal2 s 179335 -400 179391 240 0 FreeSans 6507 90 0 0 la_oenb[65]
flabel metal2 s 181108 -400 181164 240 0 FreeSans 6507 90 0 0 la_oenb[66]
flabel metal2 s 182881 -400 182937 240 0 FreeSans 6507 90 0 0 la_oenb[67]
flabel metal2 s 184654 -400 184710 240 0 FreeSans 6507 90 0 0 la_oenb[68]
flabel metal2 s 186427 -400 186483 240 0 FreeSans 6507 90 0 0 la_oenb[69]
flabel metal2 s 74728 -400 74784 240 0 FreeSans 6507 90 0 0 la_oenb[6]
flabel metal2 s 188200 -400 188256 240 0 FreeSans 6507 90 0 0 la_oenb[70]
flabel metal2 s 189973 -400 190029 240 0 FreeSans 6507 90 0 0 la_oenb[71]
flabel metal2 s 191746 -400 191802 240 0 FreeSans 6507 90 0 0 la_oenb[72]
flabel metal2 s 193519 -400 193575 240 0 FreeSans 6507 90 0 0 la_oenb[73]
flabel metal2 s 195292 -400 195348 240 0 FreeSans 6507 90 0 0 la_oenb[74]
flabel metal2 s 197065 -400 197121 240 0 FreeSans 6507 90 0 0 la_oenb[75]
flabel metal2 s 198838 -400 198894 240 0 FreeSans 6507 90 0 0 la_oenb[76]
flabel metal2 s 200611 -400 200667 240 0 FreeSans 6507 90 0 0 la_oenb[77]
flabel metal2 s 202384 -400 202440 240 0 FreeSans 6507 90 0 0 la_oenb[78]
flabel metal2 s 204157 -400 204213 240 0 FreeSans 6507 90 0 0 la_oenb[79]
flabel metal2 s 76501 -400 76557 240 0 FreeSans 6507 90 0 0 la_oenb[7]
flabel metal2 s 205930 -400 205986 240 0 FreeSans 6507 90 0 0 la_oenb[80]
flabel metal2 s 207703 -400 207759 240 0 FreeSans 6507 90 0 0 la_oenb[81]
flabel metal2 s 209476 -400 209532 240 0 FreeSans 6507 90 0 0 la_oenb[82]
flabel metal2 s 211249 -400 211305 240 0 FreeSans 6507 90 0 0 la_oenb[83]
flabel metal2 s 213022 -400 213078 240 0 FreeSans 6507 90 0 0 la_oenb[84]
flabel metal2 s 214795 -400 214851 240 0 FreeSans 6507 90 0 0 la_oenb[85]
flabel metal2 s 216568 -400 216624 240 0 FreeSans 6507 90 0 0 la_oenb[86]
flabel metal2 s 218341 -400 218397 240 0 FreeSans 6507 90 0 0 la_oenb[87]
flabel metal2 s 220114 -400 220170 240 0 FreeSans 6507 90 0 0 la_oenb[88]
flabel metal2 s 221887 -400 221943 240 0 FreeSans 6507 90 0 0 la_oenb[89]
flabel metal2 s 78274 -400 78330 240 0 FreeSans 6507 90 0 0 la_oenb[8]
flabel metal2 s 223660 -400 223716 240 0 FreeSans 6507 90 0 0 la_oenb[90]
flabel metal2 s 225433 -400 225489 240 0 FreeSans 6507 90 0 0 la_oenb[91]
flabel metal2 s 227206 -400 227262 240 0 FreeSans 6507 90 0 0 la_oenb[92]
flabel metal2 s 228979 -400 229035 240 0 FreeSans 6507 90 0 0 la_oenb[93]
flabel metal2 s 230752 -400 230808 240 0 FreeSans 6507 90 0 0 la_oenb[94]
flabel metal2 s 232525 -400 232581 240 0 FreeSans 6507 90 0 0 la_oenb[95]
flabel metal2 s 234298 -400 234354 240 0 FreeSans 6507 90 0 0 la_oenb[96]
flabel metal2 s 236071 -400 236127 240 0 FreeSans 6507 90 0 0 la_oenb[97]
flabel metal2 s 237844 -400 237900 240 0 FreeSans 6507 90 0 0 la_oenb[98]
flabel metal2 s 239617 -400 239673 240 0 FreeSans 6507 90 0 0 la_oenb[99]
flabel metal2 s 80047 -400 80103 240 0 FreeSans 6507 90 0 0 la_oenb[9]
flabel metal2 s 289852 -400 289908 240 0 FreeSans 6507 90 0 0 user_clock2
flabel metal2 s 290443 -400 290499 240 0 FreeSans 6507 90 0 0 user_irq[0]
flabel metal2 s 291034 -400 291090 240 0 FreeSans 6507 90 0 0 user_irq[1]
flabel metal2 s 291625 -400 291681 240 0 FreeSans 6507 90 0 0 user_irq[2]
flabel metal3 s 291170 319892 292400 322292 0 FreeSans 6507 0 0 0 vccd1
flabel metal3 s 291170 314892 292400 317292 0 FreeSans 6507 0 0 0 vccd1
flabel metal3 s 0 321921 830 324321 0 FreeSans 6507 0 0 0 vccd2
flabel metal3 s 0 316921 830 319321 0 FreeSans 6507 0 0 0 vccd2
flabel metal3 s 291170 270281 292400 272681 0 FreeSans 6507 0 0 0 vdda1
flabel metal3 s 291170 275281 292400 277681 0 FreeSans 6507 0 0 0 vdda1
flabel metal3 s 291170 117615 292400 120015 0 FreeSans 6507 0 0 0 vdda1
flabel metal3 s 291170 112615 292400 115015 0 FreeSans 6507 0 0 0 vdda1
flabel metal3 s 0 102444 830 104844 0 FreeSans 6507 0 0 0 vdda2
flabel metal3 s 0 107444 830 109844 0 FreeSans 6507 0 0 0 vdda2
flabel metal3 s 260297 351170 262697 352400 0 FreeSans 11166 180 0 0 vssa1
flabel metal3 s 255297 351170 257697 352400 0 FreeSans 11166 180 0 0 vssa1
flabel metal3 s 291170 73415 292400 75815 0 FreeSans 6507 0 0 0 vssa1
flabel metal3 s 291170 68415 292400 70815 0 FreeSans 6507 0 0 0 vssa1
flabel metal3 s 0 279721 830 282121 0 FreeSans 6507 0 0 0 vssa2
flabel metal3 s 0 274721 830 277121 0 FreeSans 6507 0 0 0 vssa2
flabel metal3 s 291170 95715 292400 98115 0 FreeSans 6507 0 0 0 vssd1
flabel metal3 s 291170 90715 292400 93115 0 FreeSans 6507 0 0 0 vssd1
flabel metal3 s 0 86444 830 88844 0 FreeSans 6507 0 0 0 vssd2
flabel metal3 s 0 81444 830 83844 0 FreeSans 6507 0 0 0 vssd2
flabel metal2 s 262 -400 318 240 0 FreeSans 6507 90 0 0 wb_clk_i
flabel metal2 s 853 -400 909 240 0 FreeSans 6507 90 0 0 wb_rst_i
flabel metal2 s 1444 -400 1500 240 0 FreeSans 6507 90 0 0 wbs_ack_o
flabel metal2 s 3808 -400 3864 240 0 FreeSans 6507 90 0 0 wbs_adr_i[0]
flabel metal2 s 23902 -400 23958 240 0 FreeSans 6507 90 0 0 wbs_adr_i[10]
flabel metal2 s 25675 -400 25731 240 0 FreeSans 6507 90 0 0 wbs_adr_i[11]
flabel metal2 s 27448 -400 27504 240 0 FreeSans 6507 90 0 0 wbs_adr_i[12]
flabel metal2 s 29221 -400 29277 240 0 FreeSans 6507 90 0 0 wbs_adr_i[13]
flabel metal2 s 30994 -400 31050 240 0 FreeSans 6507 90 0 0 wbs_adr_i[14]
flabel metal2 s 32767 -400 32823 240 0 FreeSans 6507 90 0 0 wbs_adr_i[15]
flabel metal2 s 34540 -400 34596 240 0 FreeSans 6507 90 0 0 wbs_adr_i[16]
flabel metal2 s 36313 -400 36369 240 0 FreeSans 6507 90 0 0 wbs_adr_i[17]
flabel metal2 s 38086 -400 38142 240 0 FreeSans 6507 90 0 0 wbs_adr_i[18]
flabel metal2 s 39859 -400 39915 240 0 FreeSans 6507 90 0 0 wbs_adr_i[19]
flabel metal2 s 6172 -400 6228 240 0 FreeSans 6507 90 0 0 wbs_adr_i[1]
flabel metal2 s 41632 -400 41688 240 0 FreeSans 6507 90 0 0 wbs_adr_i[20]
flabel metal2 s 43405 -400 43461 240 0 FreeSans 6507 90 0 0 wbs_adr_i[21]
flabel metal2 s 45178 -400 45234 240 0 FreeSans 6507 90 0 0 wbs_adr_i[22]
flabel metal2 s 46951 -400 47007 240 0 FreeSans 6507 90 0 0 wbs_adr_i[23]
flabel metal2 s 48724 -400 48780 240 0 FreeSans 6507 90 0 0 wbs_adr_i[24]
flabel metal2 s 50497 -400 50553 240 0 FreeSans 6507 90 0 0 wbs_adr_i[25]
flabel metal2 s 52270 -400 52326 240 0 FreeSans 6507 90 0 0 wbs_adr_i[26]
flabel metal2 s 54043 -400 54099 240 0 FreeSans 6507 90 0 0 wbs_adr_i[27]
flabel metal2 s 55816 -400 55872 240 0 FreeSans 6507 90 0 0 wbs_adr_i[28]
flabel metal2 s 57589 -400 57645 240 0 FreeSans 6507 90 0 0 wbs_adr_i[29]
flabel metal2 s 8536 -400 8592 240 0 FreeSans 6507 90 0 0 wbs_adr_i[2]
flabel metal2 s 59362 -400 59418 240 0 FreeSans 6507 90 0 0 wbs_adr_i[30]
flabel metal2 s 61135 -400 61191 240 0 FreeSans 6507 90 0 0 wbs_adr_i[31]
flabel metal2 s 10900 -400 10956 240 0 FreeSans 6507 90 0 0 wbs_adr_i[3]
flabel metal2 s 13264 -400 13320 240 0 FreeSans 6507 90 0 0 wbs_adr_i[4]
flabel metal2 s 15037 -400 15093 240 0 FreeSans 6507 90 0 0 wbs_adr_i[5]
flabel metal2 s 16810 -400 16866 240 0 FreeSans 6507 90 0 0 wbs_adr_i[6]
flabel metal2 s 18583 -400 18639 240 0 FreeSans 6507 90 0 0 wbs_adr_i[7]
flabel metal2 s 20356 -400 20412 240 0 FreeSans 6507 90 0 0 wbs_adr_i[8]
flabel metal2 s 22129 -400 22185 240 0 FreeSans 6507 90 0 0 wbs_adr_i[9]
flabel metal2 s 2035 -400 2091 240 0 FreeSans 6507 90 0 0 wbs_cyc_i
flabel metal2 s 4399 -400 4455 240 0 FreeSans 6507 90 0 0 wbs_dat_i[0]
flabel metal2 s 24493 -400 24549 240 0 FreeSans 6507 90 0 0 wbs_dat_i[10]
flabel metal2 s 26266 -400 26322 240 0 FreeSans 6507 90 0 0 wbs_dat_i[11]
flabel metal2 s 28039 -400 28095 240 0 FreeSans 6507 90 0 0 wbs_dat_i[12]
flabel metal2 s 29812 -400 29868 240 0 FreeSans 6507 90 0 0 wbs_dat_i[13]
flabel metal2 s 31585 -400 31641 240 0 FreeSans 6507 90 0 0 wbs_dat_i[14]
flabel metal2 s 33358 -400 33414 240 0 FreeSans 6507 90 0 0 wbs_dat_i[15]
flabel metal2 s 35131 -400 35187 240 0 FreeSans 6507 90 0 0 wbs_dat_i[16]
flabel metal2 s 36904 -400 36960 240 0 FreeSans 6507 90 0 0 wbs_dat_i[17]
flabel metal2 s 38677 -400 38733 240 0 FreeSans 6507 90 0 0 wbs_dat_i[18]
flabel metal2 s 40450 -400 40506 240 0 FreeSans 6507 90 0 0 wbs_dat_i[19]
flabel metal2 s 6763 -400 6819 240 0 FreeSans 6507 90 0 0 wbs_dat_i[1]
flabel metal2 s 42223 -400 42279 240 0 FreeSans 6507 90 0 0 wbs_dat_i[20]
flabel metal2 s 43996 -400 44052 240 0 FreeSans 6507 90 0 0 wbs_dat_i[21]
flabel metal2 s 45769 -400 45825 240 0 FreeSans 6507 90 0 0 wbs_dat_i[22]
flabel metal2 s 47542 -400 47598 240 0 FreeSans 6507 90 0 0 wbs_dat_i[23]
flabel metal2 s 49315 -400 49371 240 0 FreeSans 6507 90 0 0 wbs_dat_i[24]
flabel metal2 s 51088 -400 51144 240 0 FreeSans 6507 90 0 0 wbs_dat_i[25]
flabel metal2 s 52861 -400 52917 240 0 FreeSans 6507 90 0 0 wbs_dat_i[26]
flabel metal2 s 54634 -400 54690 240 0 FreeSans 6507 90 0 0 wbs_dat_i[27]
flabel metal2 s 56407 -400 56463 240 0 FreeSans 6507 90 0 0 wbs_dat_i[28]
flabel metal2 s 58180 -400 58236 240 0 FreeSans 6507 90 0 0 wbs_dat_i[29]
flabel metal2 s 9127 -400 9183 240 0 FreeSans 6507 90 0 0 wbs_dat_i[2]
flabel metal2 s 59953 -400 60009 240 0 FreeSans 6507 90 0 0 wbs_dat_i[30]
flabel metal2 s 61726 -400 61782 240 0 FreeSans 6507 90 0 0 wbs_dat_i[31]
flabel metal2 s 11491 -400 11547 240 0 FreeSans 6507 90 0 0 wbs_dat_i[3]
flabel metal2 s 13855 -400 13911 240 0 FreeSans 6507 90 0 0 wbs_dat_i[4]
flabel metal2 s 15628 -400 15684 240 0 FreeSans 6507 90 0 0 wbs_dat_i[5]
flabel metal2 s 17401 -400 17457 240 0 FreeSans 6507 90 0 0 wbs_dat_i[6]
flabel metal2 s 19174 -400 19230 240 0 FreeSans 6507 90 0 0 wbs_dat_i[7]
flabel metal2 s 20947 -400 21003 240 0 FreeSans 6507 90 0 0 wbs_dat_i[8]
flabel metal2 s 22720 -400 22776 240 0 FreeSans 6507 90 0 0 wbs_dat_i[9]
flabel metal2 s 4990 -400 5046 240 0 FreeSans 6507 90 0 0 wbs_dat_o[0]
flabel metal2 s 25084 -400 25140 240 0 FreeSans 6507 90 0 0 wbs_dat_o[10]
flabel metal2 s 26857 -400 26913 240 0 FreeSans 6507 90 0 0 wbs_dat_o[11]
flabel metal2 s 28630 -400 28686 240 0 FreeSans 6507 90 0 0 wbs_dat_o[12]
flabel metal2 s 30403 -400 30459 240 0 FreeSans 6507 90 0 0 wbs_dat_o[13]
flabel metal2 s 32176 -400 32232 240 0 FreeSans 6507 90 0 0 wbs_dat_o[14]
flabel metal2 s 33949 -400 34005 240 0 FreeSans 6507 90 0 0 wbs_dat_o[15]
flabel metal2 s 35722 -400 35778 240 0 FreeSans 6507 90 0 0 wbs_dat_o[16]
flabel metal2 s 37495 -400 37551 240 0 FreeSans 6507 90 0 0 wbs_dat_o[17]
flabel metal2 s 39268 -400 39324 240 0 FreeSans 6507 90 0 0 wbs_dat_o[18]
flabel metal2 s 41041 -400 41097 240 0 FreeSans 6507 90 0 0 wbs_dat_o[19]
flabel metal2 s 7354 -400 7410 240 0 FreeSans 6507 90 0 0 wbs_dat_o[1]
flabel metal2 s 42814 -400 42870 240 0 FreeSans 6507 90 0 0 wbs_dat_o[20]
flabel metal2 s 44587 -400 44643 240 0 FreeSans 6507 90 0 0 wbs_dat_o[21]
flabel metal2 s 46360 -400 46416 240 0 FreeSans 6507 90 0 0 wbs_dat_o[22]
flabel metal2 s 48133 -400 48189 240 0 FreeSans 6507 90 0 0 wbs_dat_o[23]
flabel metal2 s 49906 -400 49962 240 0 FreeSans 6507 90 0 0 wbs_dat_o[24]
flabel metal2 s 51679 -400 51735 240 0 FreeSans 6507 90 0 0 wbs_dat_o[25]
flabel metal2 s 53452 -400 53508 240 0 FreeSans 6507 90 0 0 wbs_dat_o[26]
flabel metal2 s 55225 -400 55281 240 0 FreeSans 6507 90 0 0 wbs_dat_o[27]
flabel metal2 s 56998 -400 57054 240 0 FreeSans 6507 90 0 0 wbs_dat_o[28]
flabel metal2 s 58771 -400 58827 240 0 FreeSans 6507 90 0 0 wbs_dat_o[29]
flabel metal2 s 9718 -400 9774 240 0 FreeSans 6507 90 0 0 wbs_dat_o[2]
flabel metal2 s 60544 -400 60600 240 0 FreeSans 6507 90 0 0 wbs_dat_o[30]
flabel metal2 s 62317 -400 62373 240 0 FreeSans 6507 90 0 0 wbs_dat_o[31]
flabel metal2 s 12082 -400 12138 240 0 FreeSans 6507 90 0 0 wbs_dat_o[3]
flabel metal2 s 14446 -400 14502 240 0 FreeSans 6507 90 0 0 wbs_dat_o[4]
flabel metal2 s 16219 -400 16275 240 0 FreeSans 6507 90 0 0 wbs_dat_o[5]
flabel metal2 s 17992 -400 18048 240 0 FreeSans 6507 90 0 0 wbs_dat_o[6]
flabel metal2 s 19765 -400 19821 240 0 FreeSans 6507 90 0 0 wbs_dat_o[7]
flabel metal2 s 21538 -400 21594 240 0 FreeSans 6507 90 0 0 wbs_dat_o[8]
flabel metal2 s 23311 -400 23367 240 0 FreeSans 6507 90 0 0 wbs_dat_o[9]
flabel metal2 s 5581 -400 5637 240 0 FreeSans 6507 90 0 0 wbs_sel_i[0]
flabel metal2 s 7945 -400 8001 240 0 FreeSans 6507 90 0 0 wbs_sel_i[1]
flabel metal2 s 10309 -400 10365 240 0 FreeSans 6507 90 0 0 wbs_sel_i[2]
flabel metal2 s 12673 -400 12729 240 0 FreeSans 6507 90 0 0 wbs_sel_i[3]
flabel metal2 s 2626 -400 2682 240 0 FreeSans 6507 90 0 0 wbs_stb_i
flabel metal2 s 3217 -400 3273 240 0 FreeSans 6507 90 0 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
