magic
tech sky130A
timestamp 1635362061
<< pwell >>
rect 308 -775 419 -732
<< nmos >>
rect 56 -298 156 -280
rect 56 -446 156 -428
rect 56 -612 156 -594
rect 54 -765 154 -747
rect 53 -919 153 -901
<< ndiff >>
rect 56 -248 156 -235
rect 56 -266 98 -248
rect 116 -266 156 -248
rect 56 -280 156 -266
rect 56 -312 156 -298
rect 56 -330 98 -312
rect 116 -330 156 -312
rect 56 -343 156 -330
rect 56 -396 156 -383
rect 56 -414 98 -396
rect 116 -414 156 -396
rect 56 -428 156 -414
rect 56 -460 156 -446
rect 56 -478 98 -460
rect 116 -478 156 -460
rect 56 -491 156 -478
rect 56 -562 156 -549
rect 56 -580 98 -562
rect 116 -580 156 -562
rect 56 -594 156 -580
rect 56 -626 156 -612
rect 56 -644 98 -626
rect 116 -644 156 -626
rect 56 -657 156 -644
rect 54 -715 154 -702
rect 54 -733 96 -715
rect 114 -733 154 -715
rect 54 -747 154 -733
rect 54 -779 154 -765
rect 54 -797 96 -779
rect 114 -797 154 -779
rect 54 -810 154 -797
rect 53 -869 153 -856
rect 53 -887 95 -869
rect 113 -887 153 -869
rect 53 -901 153 -887
rect 53 -933 153 -919
rect 53 -951 95 -933
rect 113 -951 153 -933
rect 53 -964 153 -951
<< ndiffc >>
rect 98 -266 116 -248
rect 98 -330 116 -312
rect 98 -414 116 -396
rect 98 -478 116 -460
rect 98 -580 116 -562
rect 98 -644 116 -626
rect 96 -733 114 -715
rect 96 -797 114 -779
rect 95 -887 113 -869
rect 95 -951 113 -933
<< psubdiff >>
rect -752 3822 -601 3831
rect -752 3781 -663 3822
rect -618 3781 -601 3822
rect -752 3772 -601 3781
rect -744 3771 -601 3772
rect 308 -745 419 -732
rect 308 -763 361 -745
rect 379 -763 419 -745
rect 308 -775 419 -763
<< psubdiffcont >>
rect -663 3781 -618 3822
rect 361 -763 379 -745
<< poly >>
rect -3 -280 31 -272
rect -3 -298 5 -280
rect 23 -298 56 -280
rect 156 -298 181 -280
rect -3 -306 31 -298
rect -3 -428 31 -420
rect -3 -446 5 -428
rect 23 -446 56 -428
rect 156 -446 181 -428
rect -3 -454 31 -446
rect -3 -594 31 -586
rect -3 -612 5 -594
rect 23 -612 56 -594
rect 156 -612 181 -594
rect -3 -620 31 -612
rect -5 -747 29 -739
rect -5 -765 3 -747
rect 21 -765 54 -747
rect 154 -765 179 -747
rect -5 -773 29 -765
rect -6 -901 28 -893
rect -6 -919 2 -901
rect 20 -919 53 -901
rect 153 -919 178 -901
rect -6 -927 28 -919
<< polycont >>
rect 5 -298 23 -280
rect 5 -446 23 -428
rect 5 -612 23 -594
rect 3 -765 21 -747
rect 2 -919 20 -901
<< locali >>
rect -4380 4217 -4324 4221
rect -4380 4171 -4374 4217
rect -4332 4171 -4324 4217
rect -4380 4114 -4324 4171
rect -4379 4087 -4324 4114
rect -1824 4202 -1768 4206
rect -1824 4156 -1818 4202
rect -1776 4156 -1768 4202
rect -1824 4099 -1768 4156
rect -4379 4078 -4322 4087
rect -4383 3997 -4322 4078
rect -1823 4072 -1768 4099
rect -1823 4063 -1766 4072
rect -4383 3853 -4320 3997
rect -1827 3982 -1766 4063
rect -4383 3847 -4315 3853
rect -4395 3812 -4312 3847
rect -1827 3812 -1764 3982
rect -766 3828 -599 3842
rect -4396 3807 -4312 3812
rect -4396 1353 -4309 3807
rect -1807 2650 -1783 3812
rect -766 3777 -738 3828
rect -688 3822 -599 3828
rect -688 3781 -663 3822
rect -618 3781 -599 3822
rect -688 3777 -599 3781
rect -766 3766 -599 3777
rect -747 3764 -610 3766
rect 2636 2688 2692 2692
rect -1807 2626 -34 2650
rect -4396 1325 -211 1353
rect -239 -390 -211 1325
rect -58 -180 -34 2626
rect 2636 2642 2642 2688
rect 2684 2642 2692 2688
rect 2636 2585 2692 2642
rect 2637 2558 2692 2585
rect 2637 2549 2694 2558
rect 2633 2380 2694 2549
rect 736 2339 2694 2380
rect -55 -206 -37 -180
rect -153 -226 -37 -206
rect -153 -254 -124 -226
rect -96 -254 -37 -226
rect -153 -281 -37 -254
rect -55 -346 -37 -281
rect -3 -248 300 -240
rect -3 -266 98 -248
rect 116 -266 300 -248
rect -3 -274 300 -266
rect -3 -280 31 -274
rect -3 -298 5 -280
rect 23 -298 31 -280
rect -3 -306 31 -298
rect 90 -312 124 -304
rect 90 -330 98 -312
rect 116 -330 124 -312
rect 90 -346 124 -330
rect -55 -368 124 -346
rect -74 -390 124 -388
rect -239 -396 124 -390
rect -239 -414 98 -396
rect 116 -414 124 -396
rect -239 -418 124 -414
rect -97 -420 124 -418
rect -97 -664 -74 -420
rect -3 -422 124 -420
rect -3 -428 31 -422
rect -3 -446 5 -428
rect 23 -446 31 -428
rect -3 -454 31 -446
rect 90 -460 124 -452
rect 90 -478 98 -460
rect 116 -478 124 -460
rect 90 -495 124 -478
rect 189 -495 209 -274
rect 270 -301 300 -274
rect 270 -346 302 -301
rect 736 -332 777 2339
rect 13729 419 14130 420
rect 13600 414 14130 419
rect 13597 412 14130 414
rect 13529 410 14130 412
rect 13395 402 14130 410
rect 13395 360 13399 402
rect 13445 360 14130 402
rect 13395 355 14130 360
rect 13395 354 13502 355
rect 13538 351 13778 355
rect 90 -527 209 -495
rect 273 -476 302 -346
rect 273 -523 575 -476
rect 544 -525 575 -523
rect 738 -525 777 -332
rect 124 -554 209 -553
rect -3 -560 209 -554
rect -3 -561 291 -560
rect 544 -561 777 -525
rect -3 -562 298 -561
rect -3 -580 98 -562
rect 116 -580 298 -562
rect -3 -588 298 -580
rect -3 -594 31 -588
rect -3 -612 5 -594
rect 23 -612 31 -594
rect -3 -620 31 -612
rect 192 -589 298 -588
rect 90 -626 124 -618
rect 90 -644 98 -626
rect 116 -644 124 -626
rect 90 -664 124 -644
rect -97 -688 124 -664
rect -226 -715 122 -707
rect -226 -733 96 -715
rect 114 -733 122 -715
rect -226 -739 122 -733
rect -226 -981 -194 -739
rect -5 -741 122 -739
rect -5 -747 29 -741
rect -5 -765 3 -747
rect 21 -765 29 -747
rect -5 -773 29 -765
rect 88 -779 122 -771
rect 88 -797 96 -779
rect 114 -797 122 -779
rect 88 -822 122 -797
rect 192 -822 209 -589
rect 248 -636 298 -589
rect 14089 -636 14130 355
rect 248 -677 14130 -636
rect 353 -745 387 -737
rect 353 -763 361 -745
rect 379 -763 387 -745
rect 353 -771 387 -763
rect -134 -858 -46 -838
rect 88 -839 209 -822
rect -134 -886 -105 -858
rect -77 -861 -46 -858
rect -77 -869 121 -861
rect -77 -886 95 -869
rect -134 -887 95 -886
rect 113 -887 121 -869
rect -134 -893 121 -887
rect -134 -913 -46 -893
rect -6 -895 121 -893
rect -6 -901 28 -895
rect -6 -919 2 -901
rect 20 -919 28 -901
rect -6 -927 28 -919
rect 87 -933 121 -925
rect 87 -951 95 -933
rect 113 -951 121 -933
rect 87 -977 121 -951
rect -39 -981 420 -977
rect -226 -1013 420 -981
rect -39 -1017 420 -1013
rect -29 -3075 55 -3073
rect -163 -3082 55 -3075
rect 380 -3082 420 -1017
rect -163 -3083 420 -3082
rect -163 -3125 -159 -3083
rect -113 -3122 420 -3083
rect -113 -3125 55 -3122
rect -163 -3130 55 -3125
rect -163 -3131 -56 -3130
rect -20 -3134 55 -3130
<< viali >>
rect -4374 4171 -4332 4217
rect -1818 4156 -1776 4202
rect -738 3777 -688 3828
rect 2642 2642 2684 2688
rect -124 -254 -96 -226
rect 13399 360 13445 402
rect -105 -886 -77 -858
rect -159 -3125 -113 -3083
<< metal1 >>
rect -4380 4217 -4324 4221
rect -4380 4171 -4374 4217
rect -4332 4171 -4324 4217
rect -4380 4143 -4324 4171
rect -1824 4202 -1768 4206
rect -1824 4156 -1818 4202
rect -1776 4156 -1768 4202
rect -1824 4128 -1768 4156
rect -763 3829 -682 3842
rect -763 3776 -738 3829
rect -688 3776 -682 3829
rect -763 3764 -682 3776
rect 2636 2688 2692 2692
rect 2636 2642 2642 2688
rect 2684 2642 2692 2688
rect 2636 2614 2692 2642
rect 13395 402 13473 410
rect 13395 360 13399 402
rect 13445 360 13473 402
rect 13395 354 13473 360
rect -153 -226 -65 -206
rect -153 -254 -124 -226
rect -96 -254 -65 -226
rect -153 -281 -65 -254
rect -134 -858 -46 -838
rect -134 -886 -105 -858
rect -77 -886 -46 -858
rect -134 -913 -46 -886
rect -163 -3083 -85 -3075
rect -163 -3125 -159 -3083
rect -113 -3125 -85 -3083
rect -163 -3131 -85 -3125
<< via1 >>
rect -4374 4171 -4332 4217
rect -1818 4156 -1776 4202
rect -738 3828 -688 3829
rect -738 3777 -688 3828
rect -738 3776 -688 3777
rect 2642 2642 2684 2688
rect 13399 360 13445 402
rect -124 -254 -96 -226
rect -105 -886 -77 -858
rect -159 -3125 -113 -3083
<< metal2 >>
rect -4380 4217 -4324 4221
rect -4380 4171 -4374 4217
rect -4332 4171 -4324 4217
rect -4380 4116 -4324 4171
rect -4380 4071 -4373 4116
rect -4331 4071 -4324 4116
rect -4380 4067 -4324 4071
rect -1824 4202 -1768 4206
rect -1824 4156 -1818 4202
rect -1776 4156 -1768 4202
rect -1824 4101 -1768 4156
rect -1824 4056 -1817 4101
rect -1775 4056 -1768 4101
rect -1824 4052 -1768 4056
rect -763 3829 -682 3842
rect -763 3776 -738 3829
rect -688 3776 -682 3829
rect -763 3764 -682 3776
rect 2636 2688 2692 2692
rect 2636 2642 2642 2688
rect 2684 2642 2692 2688
rect 2636 2587 2692 2642
rect 2636 2542 2643 2587
rect 2685 2542 2692 2587
rect 2636 2538 2692 2542
rect 13395 403 13549 410
rect 13395 402 13500 403
rect 13395 360 13399 402
rect 13445 361 13500 402
rect 13545 361 13549 403
rect 13445 360 13549 361
rect 13395 354 13549 360
rect -153 -226 -65 -206
rect -153 -254 -124 -226
rect -96 -254 -65 -226
rect -153 -281 -65 -254
rect -134 -858 -46 -838
rect -134 -886 -105 -858
rect -77 -886 -46 -858
rect -134 -913 -46 -886
rect -110 -1135 -56 -913
rect -110 -1183 1399 -1135
rect -163 -3082 -9 -3075
rect -163 -3083 -58 -3082
rect -163 -3125 -159 -3083
rect -113 -3124 -58 -3083
rect -13 -3124 -9 -3082
rect -113 -3125 -9 -3124
rect -163 -3131 -9 -3125
rect 1351 -4539 1399 -1183
rect 1811 -4508 1976 -4472
rect 1811 -4539 1855 -4508
rect 1351 -4587 1855 -4539
rect 1811 -4603 1855 -4587
rect 1949 -4603 1976 -4508
rect 1811 -4649 1976 -4603
<< via2 >>
rect -4373 4071 -4331 4116
rect -1817 4056 -1775 4101
rect -738 3777 -688 3828
rect 2643 2542 2685 2587
rect 13500 361 13545 403
rect -124 -254 -96 -226
rect -58 -3124 -13 -3082
rect 1855 -4603 1949 -4508
<< metal3 >>
rect -5522 17020 -2930 17059
rect -4403 4230 -3875 14258
rect -3945 4158 -3903 4230
rect -4380 4116 -4324 4122
rect -4380 4071 -4373 4116
rect -4331 4071 -4324 4116
rect -4380 4067 -4324 4071
rect -3944 3827 -3905 4158
rect -3943 -1419 -3905 3827
rect -2969 722 -2930 17020
rect -1847 4215 -1319 14243
rect -1389 4143 -1347 4215
rect -1824 4101 -1768 4107
rect -1824 4056 -1817 4101
rect -1775 4056 -1768 4101
rect -1824 4052 -1768 4056
rect -1388 3853 -1349 4143
rect -1388 3749 -1347 3853
rect -743 3845 -683 17075
rect -743 3828 -681 3845
rect -743 3777 -738 3828
rect -688 3777 -681 3828
rect -743 3771 -681 3777
rect -744 3749 -681 3771
rect -1388 3742 -681 3749
rect -1388 3692 -685 3742
rect 2613 2701 3141 12729
rect 3071 2629 3113 2701
rect 2636 2587 2692 2593
rect 2636 2542 2643 2587
rect 2685 2542 2692 2587
rect 2636 2538 2692 2542
rect 3071 2307 3106 2629
rect 3070 1277 3106 2307
rect 13808 1277 13844 3144
rect 3070 1241 13844 1277
rect 3358 831 13386 859
rect 3358 825 13458 831
rect 13808 825 13844 1241
rect 3358 789 13844 825
rect -2969 683 -356 722
rect -395 -223 -356 683
rect 3358 331 13386 789
rect 13494 403 13549 410
rect 13494 361 13500 403
rect 13545 361 13549 403
rect 13494 354 13549 361
rect -153 -223 -65 -206
rect -395 -226 -65 -223
rect -395 -254 -124 -226
rect -96 -254 -65 -226
rect -395 -262 -65 -254
rect -177 -263 -65 -262
rect -153 -281 -65 -263
rect -133 -282 -92 -281
rect -3943 -1420 760 -1419
rect -3943 -1457 826 -1420
rect 781 -1630 826 -1457
rect 781 -1962 817 -1630
rect 16523 -1962 16559 3105
rect 781 -1998 16559 -1962
rect -10200 -2654 -172 -2626
rect -10200 -2660 -100 -2654
rect 781 -2660 817 -1998
rect -10200 -2696 817 -2660
rect -10200 -3154 -172 -2696
rect -64 -3082 -9 -3075
rect -64 -3124 -58 -3082
rect -13 -3124 -9 -3082
rect -64 -3131 -9 -3124
rect 1811 -4503 1976 -4472
rect 1811 -4508 2140 -4503
rect 1811 -4603 1855 -4508
rect 1949 -4603 2140 -4508
rect 1811 -4614 2140 -4603
rect 1811 -4649 1976 -4614
<< via3 >>
rect -4373 4071 -4331 4116
rect -1817 4056 -1775 4101
rect 2643 2542 2685 2587
rect 13500 361 13545 403
rect -58 -3124 -13 -3082
<< mimcap >>
rect -4389 4289 -3889 14244
rect -4389 4256 -4366 4289
rect -4333 4256 -3889 4289
rect -4389 4244 -3889 4256
rect -1833 4274 -1333 14229
rect -1833 4241 -1810 4274
rect -1777 4241 -1333 4274
rect -1833 4229 -1333 4241
rect 2627 2760 3127 12715
rect 2627 2727 2650 2760
rect 2683 2727 3127 2760
rect 2627 2715 3127 2727
rect 3372 401 13372 845
rect 3372 368 13327 401
rect 13360 368 13372 401
rect 3372 345 13372 368
rect -10186 -3084 -186 -2640
rect -10186 -3117 -231 -3084
rect -198 -3117 -186 -3084
rect -10186 -3140 -186 -3117
<< mimcapcontact >>
rect -4366 4256 -4333 4289
rect -1810 4241 -1777 4274
rect 2650 2727 2683 2760
rect 13327 368 13360 401
rect -231 -3117 -198 -3084
<< metal4 >>
rect -4372 4289 -4327 4298
rect -4372 4256 -4366 4289
rect -4333 4256 -4327 4289
rect -4372 4221 -4327 4256
rect -1816 4274 -1771 4283
rect -1816 4241 -1810 4274
rect -1777 4241 -1771 4274
rect -4380 4116 -4324 4221
rect -1816 4206 -1771 4241
rect -4380 4071 -4373 4116
rect -4331 4071 -4324 4116
rect -4380 4068 -4324 4071
rect -1824 4101 -1768 4206
rect -1824 4056 -1817 4101
rect -1775 4056 -1768 4101
rect -1824 4053 -1768 4056
rect 2644 2760 2689 2769
rect 2644 2727 2650 2760
rect 2683 2727 2689 2760
rect 2644 2692 2689 2727
rect 2636 2587 2692 2692
rect 2636 2542 2643 2587
rect 2685 2542 2692 2587
rect 2636 2539 2692 2542
rect 13395 407 13548 410
rect 13318 403 13548 407
rect 13318 401 13500 403
rect 13318 368 13327 401
rect 13360 368 13500 401
rect 13318 362 13500 368
rect 13395 361 13500 362
rect 13545 361 13548 403
rect 13395 354 13548 361
rect -163 -3078 -10 -3075
rect -240 -3082 -10 -3078
rect -240 -3084 -58 -3082
rect -240 -3117 -231 -3084
rect -198 -3117 -58 -3084
rect -240 -3123 -58 -3117
rect -163 -3124 -58 -3123
rect -13 -3124 -10 -3082
rect -163 -3131 -10 -3124
<< labels >>
rlabel metal3 -139 -241 -139 -241 1 io_analog[2]
rlabel via2 -715 3807 -715 3807 1 vssa1
rlabel metal2 -87 -904 -87 -904 1 vccd1
rlabel metal3 800 -1979 800 -1979 1 io_analog[0]
rlabel metal3 13823 1255 13823 1255 1 io_analog[1]
<< end >>
